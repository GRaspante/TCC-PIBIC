----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 09.04.2023 12:24:00
-- Design Name: 
-- Module Name: fpupack - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;
package fpupack is
    constant FRAC_WIDTH : integer := 18;
    constant EXP_WIDTH : integer := 8;
    constant FP_WIDTH : integer:= FRAC_WIDTH+EXP_WIDTH+1;
    constant bias : std_logic_vector(EXP_WIDTH-1 downto 0) := "01111111";
    constant int_bias : integer := 127;
    constant int_alin : integer := 255;
    constant EXP_DF : std_logic_vector(EXP_WIDTH-1 downto 0) := "10000010";
    constant bias_MAX : std_logic_vector(EXP_WIDTH-1 downto 0) := "10000110";
    constant bias_MIN : std_logic_vector(EXP_WIDTH-1 downto 0) := "01110101";
    constant EXP_ONE: std_logic_vector(EXP_WIDTH-1 downto 0):= (others => '1');
    constant EXP_INF : std_logic_vector(EXP_WIDTH-1 downto 0) := "11111111";
    constant ZERO_V : std_logic_vector(FP_WIDTH-1 downto 0) := (others => '0');
   
    constant s_one : std_logic_vector(FP_WIDTH-1 downto 0) := "001111111000000000000000000";                                                               
    constant s_ten : std_logic_vector(FP_WIDTH-1 downto 0) := "010000010010000000000000000";                      
    constant s_twn : std_logic_vector(FP_WIDTH-1 downto 0) := "010000011010000000000000000";
    constant s_hundred : std_logic_vector(FP_WIDTH-1 downto 0) := "010000101100100000000000000";                                                                   
    constant s_pi2 : std_logic_vector(FP_WIDTH-1 downto 0) := "001111111100100100001111110";
    constant s_pi : std_logic_vector(FP_WIDTH-1 downto 0) := "010000000100100100001111110";
    constant s_3pi2 : std_logic_vector(FP_WIDTH-1 downto 0) := "010000001001011011001011111";
    constant s_2pi : std_logic_vector(FP_WIDTH-1 downto 0) := "010000001100100100001111110";
    
    constant Phyp : std_logic_vector(FP_WIDTH-1 downto 0) := "001111111001101001000001111";
    constant log2e : std_logic_vector(FP_WIDTH-1 downto 0) := "001111111011100010101010001";
    constant ilog2e : std_logic_vector(FP_WIDTH-1 downto 0) := "001111110011000101110010000";
    constant d_043 : std_logic_vector(FP_WIDTH-1 downto 0) :=  "001111010011000000100000110";
   
    constant MAX_ITER_CORDIC : std_logic_vector(4 downto 0):= "01111";
    constant MAX_POLY_MACKLR : std_logic_vector(3 downto 0):= "0011";
   
    constant OneM: std_logic_vector(FRAC_WIDTH downto 0) := "1000000000000000000";
    constant Zero: std_logic_vector(FP_WIDTH-1 downto 0) := (others => '0');
    constant Inf: std_logic_vector(FP_WIDTH-1 downto 0) := "011111111000000000000000000";
    constant NaN: std_logic_vector(FP_WIDTH-1 downto 0) := "011111111100000000000000000";
    constant TSed: POSITIVE := 15;
    constant Niter: POSITIVE := 3;
    
    -- PARAMETROS DA DIMEN��O DA CAMADA CONVOLUCIONAL
    constant sampleLength : integer := 66;
    constant numberOfFilters : integer := 32;
    constant biasConvLength : integer := 32;
    
   -- ARRAYS PARA A PRIMEIRA CAMADA DE CONVOLU��O
    TYPE samples_adjust IS ARRAY ((sampleLength-1) downto 0) of std_logic_vector ((FP_WIDTH - 1) downto 0);
    TYPE filter IS ARRAY ((numberOfFilters-1) downto 0, 6 downto 0) of std_logic_vector ((FP_WIDTH-1) downto 0);
    TYPE biasConv IS ARRAY ((biasConvLength-1) downto 0) of std_logic_vector ((FP_WIDTH-1) downto 0);
    TYPE outConv IS ARRAY ((numberOfFilters-1) downto 0, 59 downto 0) of std_logic_vector ((FP_WIDTH-1) downto 0);

    -- CONSTANTES DOS FILTROS E BIAS ARMAZENADOS EM BROM DA FPGA
    constant firstConvFilter : filter := (("101111100011011000101000011","101111100010010010010000000","001111001000110100101100000","101111010101001110110011101","101111100011100101000101111","101111011011101011111110100","101111100011101010011100010"),
    ("101111100000001010110010001","001111001001111110111010100","001111000110011101100011100","001111100000010000100101011","101111011110001100000001010","001111011101010011000010100","101111001100010001001000000"),
    ("101111100100000101001100011","101111100010101011100101000","101111011111101001101100000","001110011100000100101000001","101111010010001001100001001","101111100010010111111100011","101111100011000111110100000"),
    ("101111011110010110010111001","101111010000001010100001000","101111100111100000111100100","101111100101001001011111011","101111100010011111000001000","101111011100011111100110011","101111100011011011100000111"),
    ("001111011111011100001101000","001111011000000111111111100","001111011001110011101010110","001110111000011001000100001","101111100000010110110000100","101111011001001001101100100","101111011101010110110111010"),
    ("001111000010010100011000001","101111011101100101110101101","001111001110001000111100011","101111010110110011101010110","101111011010100011011011111","001111100000011100100100000","001111010000011100101101001"),
    ("101111001000111010000111001","101111100000011001101101100","101111100100111001000101101","101111010100100000100101111","101111011001111110110100100","101111011101101001000010001","101111100010111111100111000"),
    ("101111100101011001010011010","001111010111001010000000000","101111010001111011101101010","101111010000110100110101001","001111011001001100100001100","001111100000000111100000110","001111100010101100100111110"),
    ("101111010100000010111111101","001111100010010001000111001","001111010010000111110000011","001110101000011110001000111","001111011111100001001001101","001111011101100101110101001","001111100001001000011001010"),
    ("101111100001001000001000010","101111100000001010010000000","101111011011001100010110100","001111100001010010101111100","101111001100110110101101001","001111100000100101110000100","101111010011101101111000100"),
    ("101111100000001100000001101","001111011011111011001110011","101111011001110011001101001","001111011111100000011101011","001110101100001000111101111","101111011011111000100000010","001111011100011000111110011"),
    ("101111010010100000011100110","101111011101101000000111111","001111010111101101100111000","001111100000010000000011010","001111100000001011111000110","101111011110001101110010011","001111010001101011010000110"),
    ("101111011101001101101000100","101111010000001101011010111","001110101000100001100010111","101111011111000001000000011","001111011111110000010001111","001111100010100000101101100","101111011001101111011111011"),
    ("101111100010100101101100100","101111010111111100100010000","101111100000010010100110101","001111011011110010011010100","101111011000011011110100001","101111100100010110101110111","101111011011100000001100111"),
    ("001111010001010111111110101","101111011100110000010001000","001111100010011101001000100","001111011100100011010011001","001111011000001111000001010","001111001010010100011101000","001111011111010001000001111"),
    ("101111010000001100010111000","101110110010000011000000110","101111001111010001110001111","001111010010110101011101011","101111010110010000001101001","001111010110001111001010100","001111011111011010100011010"),
    ("001111011001100010001100001","101111010001100110100110100","101111010010100001011110010","001111000011110001010000001","001111001111111100110000110","101111011101100000000100101","001111010011001110101101011"),
    ("001111100001000011010001110","001111100000000101010110110","001111011001110111001001100","001111011111000101101111000","001111100001110101000001001","001111011011111100100111010","001111011000001111011010110"),
    ("101111000010101001011011001","001111001000100000100000111","001111011010011001011011010","001110111110100011001010010","001111010100100010101001001","001111011111111010010110100","101111100010010101111100110"),
    ("101111100101100011011001000","101111010100001110100101101","001111010100010001101010100","101111011001101011111101000","001111011000011011110010000","101111010011011011010001001","101111011011001000100100011"),
    ("101111001000011001100100000","101111010011101100010111111","001111001010001100101101110","101111010110111111011101000","101111011101101010110000110","101111100101111100100010111","101111100100111001110000000"),
    ("101111010110100001110000110","001111011001101010111011010","101111001011111001011001001","101110110010000010001001100","101111100011101011011100001","001111001110010000011111000","101111100011100100101010000"),
    ("001111100000010111101001000","001111010100110101000000000","001111011011010110010111010","101111011111111000000001000","101111011101111111011101110","101111000101100001001110110","101111011110101110110110001"),
    ("001111000101111100100001101","101111100001110000110000011","101111100010000010000011001","101111100101101001101110101","001110101011010001011100001","101111010011110101010000101","101111011001000011101101011"),
    ("101111011111111010111101100","001111011011101000000000001","001111011110100010101010111","001111100000100010001010001","101111011010000101001101111","001111011010110110110110111","101111100000011100001001101"),
    ("101111011000000001001100011","101111011010011001110111001","001111011110000100011010000","001111010101100100000100001","101111011000101001001100100","101111001001101101110111101","001111001011100100000011010"),
    ("001111100001111110011111100","101111011010101110000100001","101111100000111011011001101","101111011011001110101010111","001111100000110100101110001","101111100000111100000110100","001111011110000101101110001"),
    ("101111010001100001111001000","001111100000101111101101000","001111011101111001100110011","001111011100001111010110110","101111010001001010110111010","001111010101111111110000100","001111011011111111110100011"),
    ("101111100001111101011010001","101111100000010110110111010","101111100000110100010001101","001111011111110100001000101","001111100010110100011011010","001111100001111001010001100","001111100001010011110100010"),
    ("101111100001101101101011101","001111011100010011010110000","101111011101100111011111010","101111011000101011100001010","001111011000000000001000011","001111010110010000101111010","001111010000111100000011011"),
    ("101111011101000110010011011","101111010000001100101101011","001111010101001011010010100","101111001100000000100001011","001111011001100010100101010","101111010000101100010110010","101111010001100111111101101"),
    ("101111011001110111010101100","101111011011110100100101010","101111010011110010110111111","101111100000111110111001111","001111011100001101101110001","001111001110001111110001001","101111011010110011110000011"));


    constant firstConvBias : biasConv := ("001110111001101011101101110","001111010011110000111000001","101110101011110110110110110","101111000000001101110110101","001111010001010010001110000","001111010110101100110011010","101110110100110010001101101","001110111100001111010100010","101111001010110000000100000","001111010110011001001100010","001111010010000000010000110","001111010000010000011011010","001111010011011011000111000","101110110101001001100010100","001111010001000011110001001","001111010101000010010111001","001111010001000111110100111","101111001010101010101101110","001111000000000111000110111","101111001000111101011101011","101110111011000100000010001","001111010010100010100001111","001111010110101101010010000","101110111000100010111111010","001111010011110111010010011","001111010101100010101100110","001111010010001010111011100","101111001001001011101101010","001111001010101110100001011","001111010010100110101100011","001111000011110011101010101","001111010100110111111010111");



end fpupack;

package body fpupack is
end fpupack;