----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 09.04.2023 12:24:00
-- Design Name: 
-- Module Name: fpupack - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;
package fpupack is
    constant FRAC_WIDTH : integer := 18;
    constant EXP_WIDTH : integer := 8;
    constant FP_WIDTH : integer:= FRAC_WIDTH+EXP_WIDTH+1;
    constant bias : std_logic_vector(EXP_WIDTH-1 downto 0) := "01111111";
    constant int_bias : integer := 127;
    constant int_alin : integer := 255;
    constant EXP_DF : std_logic_vector(EXP_WIDTH-1 downto 0) := "10000010";
    constant bias_MAX : std_logic_vector(EXP_WIDTH-1 downto 0) := "10000110";
    constant bias_MIN : std_logic_vector(EXP_WIDTH-1 downto 0) := "01110101";
    constant EXP_ONE: std_logic_vector(EXP_WIDTH-1 downto 0):= (others => '1');
    constant EXP_INF : std_logic_vector(EXP_WIDTH-1 downto 0) := "11111111";
    constant ZERO_V : std_logic_vector(FP_WIDTH-1 downto 0) := (others => '0');
   
    constant s_one : std_logic_vector(FP_WIDTH-1 downto 0) := "001111111000000000000000000";                                                               
    constant s_ten : std_logic_vector(FP_WIDTH-1 downto 0) := "010000010010000000000000000";                      
    constant s_twn : std_logic_vector(FP_WIDTH-1 downto 0) := "010000011010000000000000000";
    constant s_hundred : std_logic_vector(FP_WIDTH-1 downto 0) := "010000101100100000000000000";                                                                   
    constant s_pi2 : std_logic_vector(FP_WIDTH-1 downto 0) := "001111111100100100001111110";
    constant s_pi : std_logic_vector(FP_WIDTH-1 downto 0) := "010000000100100100001111110";
    constant s_3pi2 : std_logic_vector(FP_WIDTH-1 downto 0) := "010000001001011011001011111";
    constant s_2pi : std_logic_vector(FP_WIDTH-1 downto 0) := "010000001100100100001111110";
    
    constant Phyp : std_logic_vector(FP_WIDTH-1 downto 0) := "001111111001101001000001111";
    constant log2e : std_logic_vector(FP_WIDTH-1 downto 0) := "001111111011100010101010001";
    constant ilog2e : std_logic_vector(FP_WIDTH-1 downto 0) := "001111110011000101110010000";
    constant d_043 : std_logic_vector(FP_WIDTH-1 downto 0) :=  "001111010011000000100000110";
   
    constant MAX_ITER_CORDIC : std_logic_vector(4 downto 0):= "01111";
    constant MAX_POLY_MACKLR : std_logic_vector(3 downto 0):= "0011";
   
    constant OneM: std_logic_vector(FRAC_WIDTH downto 0) := "1000000000000000000";
    constant Zero: std_logic_vector(FP_WIDTH-1 downto 0) := (others => '0');
    constant Inf: std_logic_vector(FP_WIDTH-1 downto 0) := "011111111000000000000000000";
    constant NaN: std_logic_vector(FP_WIDTH-1 downto 0) := "011111111100000000000000000";
    constant TSed: POSITIVE := 15;
    constant Niter: POSITIVE := 3;
    
    -- PARAMETROS DA DIMEN��O DA CAMADA CONVOLUCIONAL
    constant sampleLength : integer := 66;
    constant inConvs : integer := 34;
    constant inConvs2 : integer := 32;
    constant outConvs : integer := 30;
    constant numberOfFilters : integer := 32;
    constant biasConvLength : integer := 32;
    
   -- ARRAYS PARA A PRIMEIRA CAMADA DE CONVOLU��O
    TYPE samples_adjust IS ARRAY ((sampleLength-1) downto 0) of std_logic_vector ((FP_WIDTH - 1) downto 0);
    TYPE filter IS ARRAY ((numberOfFilters-1) downto 0, 6 downto 0) of std_logic_vector ((FP_WIDTH-1) downto 0);
    TYPE biasConv IS ARRAY ((biasConvLength-1) downto 0) of std_logic_vector ((FP_WIDTH-1) downto 0);
    TYPE outConv IS ARRAY ((numberOfFilters-1) downto 0, 59 downto 0) of std_logic_vector ((FP_WIDTH-1) downto 0);
    -- ARRAYS PARA A SEGUNDA CAMADA DE CONVOLU��O
    TYPE in_Conv2 IS ARRAY ((numberOfFilters-1) downto 0, (inConvs-1) downto 0) of std_logic_vector ((FP_WIDTH-1) downto 0);
    TYPE filter2 IS ARRAY ((numberOfFilters-1) downto 0, (numberOfFilters-1) downto 0, 4 downto 0) of std_logic_vector ((FP_WIDTH-1) downto 0);
    TYPE aux_filter2 IS ARRAY ((numberOfFilters-1) downto 0, 4 downto 0) of std_logic_vector ((FP_WIDTH-1) downto 0);
    TYPE out_loop IS ARRAY ((numberOfFilters-1) downto 0) of std_logic_vector ((FP_WIDTH-1) downto 0);
    TYPE out_Conv2 IS ARRAY ((numberOfFilters-1) downto 0, (outConvs-1) downto 0) of std_logic_vector ((FP_WIDTH-1) downto 0);
    -- ARRAYS PARA A TERCEIRA CAMADA DE CONVOLU��O
    TYPE in_Conv3 IS ARRAY ((numberOfFilters-1) downto 0, (inConvs2-1) downto 0) of std_logic_vector ((FP_WIDTH-1) downto 0);
    TYPE filter3 IS ARRAY ((numberOfFilters-1) downto 0, (numberOfFilters-1) downto 0, 2 downto 0) of std_logic_vector ((FP_WIDTH-1) downto 0);
    TYPE aux_filter3 IS ARRAY ((numberOfFilters-1) downto 0, 2 downto 0) of std_logic_vector ((FP_WIDTH-1) downto 0);

  
    -- CONSTANTES DOS FILTROS E BIAS ARMAZENADOS EM BROM DA FPGA
   
    constant thirdConvBias : biasConv := ("001111011000111011111010111","001111001001010011110111000","101111001100001111011011001","001111000000001000111111011","101111001101011101110001010","101110011100001011010100011","001111010010111000101110001","001111001011101100111001011","101111001101010111111111101","101111000000010011010011111","001111001010100111000111101","101111010111011000001010110","101110111100110111010000001","001111010001011100010111010","001111001001010100101101010","101110111111001110010110000","101110110010010001111110110","001111010111001011011001000","001110110000101100101110101","001111001111001111001010010","001110111100111000111101001","001111010000100001101011110","001111001000101001101001100","001111000111101010011000101","101111001010000011100011111","101110111110011110001111000","001111001100110110100001011","001111001001101100111101101","001111001110110110101001001","001110111011100010110101011","101111000110111100101111000","001111010010101000110001011");

constant thirdConvfilter : filter3 :=((("101111010111010000110100100","001111011100101111011011011","101111001101111011000111011"),
("101111010110001101000111000","101111100000000001101110010","101111100000001000111000101"),
("101111100001010101100110111","001111100010111100001101011","101111011010110001001101111"),
("101111100011100110000100100","101111011110001010010010010","001111010001110000100111110"),
("101111011000011110101101111","001111011001001000111100000","001111100011000110100100001"),
("101111100000100100100110010","101111011011011101111011100","001111011001010110101011111"),
("101111000100000100101100100","001111100000100110110011001","001111100100010010001111110"),
("001111100000001101001000010","101111011100011010001011000","001111100000111000010101110"),
("101111011100011100011000101","001111100001101001000000000","001111001000110011111111111"),
("101111011110111100010110000","001111100101101100110000111","001111100100001111110101111"),
("001111011110100000101111001","101111001010010101100110011","001110111101101001101010100"),
("101111001110101000111101010","101111011010110011111010010","001111010110000111011000101"),
("001111100010111110010111101","001111011110011111100001111","001111100000100100001010010"),
("101111001111110001010011110","001111010111011000001000000","101111100001101111101101110"),
("001111010100010001011000010","001111010001110001010010101","001111011110100110111111101"),
("001111001010011011010100101","001111011101001011100110100","101111010011100100010111101"),
("001111011100000010110010001","101111010110001100100000000","001111000010100000111101110"),
("101111010101001110111100010","001111100010010100000100001","101111010010001110101010100"),
("001111100010101111010011101","001111011010111111010010110","101111001101100110111011111"),
("101111010000000000111000001","001110111000110110111101000","001111011111110101000101001"),
("001111100010110111001011010","001111010101101001111111100","001111100100011010010110000"),
("101111011100010110111010001","001111010111001001100010000","001111100000010001111001101"),
("101111011000100010110011000","101111010100100010000110111","101111100000000001001000010"),
("101111100001010001100110010","001111100000001100111111011","101111011001110010111111000"),
("001111100010000111100000101","001111100000101110110001100","101111001110101101010000011"),
("001111010000101001101001101","001111010111001110110001010","101111001110001000100111101"),
("001111100001011010000101101","101111011001010100010010000","001111100001011001001001001"),
("001111011111011111011101101","001111011011100000000010011","001111011101000100000101100"),
("001111100101000011110001100","001111011011110111000111001","101111001011000110000000111"),
("001111011110000001110111111","001111010010100011101011101","101111100011101110110010111"),
("001111011010101010110010110","101111010011101001101111000","001111010001101011011100111"),
("101111100000010011111011011","101111100110110110101110101","101111011101110000010110111")),
(("001111011011101101011001011","001111100100011110000110001","101111100001101101110001010"),
("101111011101011010111111111","101111100010000000010011101","101111010011010110111010001"),
("001111100101001010010100101","001111011101100100010110010","101111011010010100100010010"),
("101111011110110010110001001","001111011101100000011110101","101111010111011011001111111"),
("101111011000101000001011100","001111100001001100100001000","001111011011111010001011010"),
("001111001110101111000010110","001111011110010110100101111","101111011010011011011110100"),
("001111011101111111110001000","001111010000101110001110011","101111010011110101000100001"),
("101111100000011100001010101","101111011010101000100011101","001111011101001011011001001"),
("101111011010010001101010000","101111010100001100011000010","101111011001100101001111010"),
("101111100101110011010111011","101110111110110000011100000","001111000111011100010010011"),
("101111100111000011100101100","101111100100101000000111011","001111011110110001000011010"),
("001111011100001101101101110","001110110010011001100001101","101111001101100101111100110"),
("001111100110110001000111010","101111010010100010011100110","101111100001000111010010000"),
("101111011111111001111101011","101111011001101110011010110","001111001010010111010011001"),
("101111011000100010111001000","101110111010011010010000100","101111001111000001010011000"),
("101111100111010000100011111","101111100010101110011110100","001111011001110111111000000"),
("001111100100101100001111000","001111100000100111111000101","101111100000001101011101010"),
("101111100010100101010000011","001111010000101001000101000","001110110000001001000001100"),
("001111011000110010100010100","001111001101010111100000111","101111011000100111101000011"),
("101111100001101100110001000","001111011011000110101100000","101111010000101000000111111"),
("101111010011101100010011110","001111100011110111111111100","001110111111010001000100110"),
("101111010110110100010000000","101111100011100101000111111","101111010010001010101101000"),
("101111010101011100000101110","001111100001100001101011101","101111100101101111000110110"),
("001111001001110000100001010","001111011010101110101000110","101111011001000000100100110"),
("101111011010001101011000000","101111100000011010111000000","001111011001110100011010111"),
("101111010011100100111100000","001111100001001101010010110","001111100001010011000110111"),
("001111011111001011110100101","001111010100010001010110001","101111100010001101111011001"),
("101111011000001000111000111","101111100010110111000110011","001111011111011100010011001"),
("001111011101101001010000111","101111000011101101110110000","101111011000101111101010100"),
("101111100000000010010010101","001111011000010101110000001","101111101001110101010000111"),
("101111011111100001010111001","101111011100111011111010111","001111100010001011001101000"),
("101111011101011001001000101","101111011010100010000101000","001111100000110010110011010")),
(("101111100000000011001100011","101111011111001110111111111","001111010111110101011010010"),
("001111011111000101010010010","001111100010100100101111110","101111010010011001111100000"),
("001111001011011010010011101","001111100111010011100110111","001111011001100001111110100"),
("101111011010111100111111001","101111011001011010101110010","001111100000111101001110111"),
("001111011010101101101101101","101111100000111101110001010","101111100100111000111100001"),
("001111100011011010010101010","101111011101001110111000110","001111011100000000010100011"),
("101111010101001111001001001","101111100000001010111010001","101111010010000110111010001"),
("001111011101001100000001010","101111010001101101001010100","001111011111100101111011111"),
("101111010000011001001100111","001111100000110000000110111","101111100001010110101001100"),
("101111011111011000100011101","101111100010010001101101110","101111001010010001010110010"),
("101111011101100101110111010","001111011110001100101010101","101111011010011100010111010"),
("101111100100000011100010110","001111100001001111100111110","101111001010000010000101111"),
("101111001101100011010100110","001111010011110110111101100","001110111101010101100011110"),
("101111011101111011011011110","001111100010010000100110001","001111011111010110011111100"),
("001111010101000100111110010","101111100000100110100000100","001111001010010111100101010"),
("001111010000100011000101110","101110111001000100011111101","001110111110100000001000000"),
("001111100010111111111100011","101111010100101001010110001","001111100001101100111100001"),
("101111011110011100000001000","101111000101011000100000100","101111011000111010011001101"),
("101111100001101000110000110","101111011101001001011011101","001111010110000110001110001"),
("101111011010001000011110110","101111011010010010010100000","001111001110010110100100100"),
("101111100001111001101010100","101111011001111000101100001","001111100010111011100010011"),
("101111010011000010100010111","001111011000001010111000010","101111100000101100111010000"),
("001111010111110001100111000","101111011100100000011101010","101111011010001110100011011"),
("101111010101101001101011010","101110110100001011111101101","101111100001000001010011110"),
("101111100001111001100001010","101111001101100011101101111","101111100000100001010100100"),
("101111011111101111010110010","001111011101110010010010010","001111011111100000011001001"),
("001111001011000000111101011","101111010001101101001000000","001111100010010101110110100"),
("001111011001100110010000011","101111011011011111110000100","101111011101110110001110101"),
("101111100011011000001101100","001111011111011010010101101","001111100000010111111011011"),
("101111011100101101111101001","001111011010001111000101101","101111011000101111010001111"),
("001111011010110111100010101","101111100101100010000101010","101111011011001110011110000"),
("101111011001001101011010101","101111100100111101100101100","001111010011000111001010100")),
(("101110111111011111110110101","101111010111110100011110101","101111011101111011010111101"),
("101111010000101001101101111","001111010100111000010010110","101111011101000001001001000"),
("001111100000010010110011010","101111010111010000110111011","001111010111011101001111101"),
("001111011010111110010011001","001111010100101010110101110","101111011000110011001000011"),
("001111011010011110100100111","001111011100010011011110110","001111010100000101111010110"),
("001111011010110011110101000","001111011001111110000100101","001111001110111001100010010"),
("001111100001001010110110100","101111010001001101101100011","101111011000101000010110110"),
("101111011010110001001100100","001111011100001000000000000","101111011101100100010001001"),
("001111001011111101001101111","001111010000010110111011100","101111011000110101111011101"),
("101111011000010101001100101","001111010001001010111110100","101111010111000100100111001"),
("001110111000110100110101111","001111100001110001011101100","101111011100111111101010111"),
("101110110110111110011011010","101111000101011001111111001","001111011100000001001110110"),
("101111010010010000101010001","001111011110011111101101110","101111011100001111110100110"),
("101111011111000100100101101","001111100001101110101110010","101111001101011001101001001"),
("101111100100010100010100100","101111010110011101010110011","101111100000011000111001111"),
("101111010100001100000001011","001111100100011101001010000","001111001011001001000011011"),
("001111100001001111111010110","101111010100000001111011001","001111011000111101000010011"),
("101111100011001110101110101","001111011100011001110110000","001111011000101110011011110"),
("101111010000001011010101010","101110111010100001000111100","001111011110000011100101111"),
("001111001110101110110111100","101111100001100110011011010","001111001000010110010000010"),
("101111010011100000101110000","001111011110010000111001000","101111010110110001111010101"),
("101111011110101101000100100","101111011010101001011001010","101111011101010001100110011"),
("001111001010010000001101001","001111000101100000001010001","101111011011110110111101110"),
("001111100011100100101011010","001111010000101101110000010","001110111100011111111011010"),
("101111100010101110010011110","101111001001011010111001000","101111100010001011001101001"),
("001111100011100011011101100","001111011000001010111100011","101111100001111010011011010"),
("001111011111111001011010111","101111010100100110101000011","001111100000011010000010101"),
("101110111001010100110101001","001111100001010111100101101","001111100010010001101011000"),
("101111100011011110100111011","001111100000100110100001110","001111100000000100111111011"),
("001111011100100000100011110","001111011101110000101010110","101111010110111100110001110"),
("101110101001000100101001101","001111011110110001111000110","101111010110010101000101010"),
("101111011001000001101010010","001111010010011110100010111","001111011100010001100111010")),
(("001110111101110100011001100","101111011110001101000011110","101111011111100110000011001"),
("101111100001110100010111111","001110110011010101100001010","001111100011100110000001001"),
("001111011000100011000111101","101111001101110110010111001","101111100000000011111000110"),
("101110111001001001001101011","101111100011101001000001010","101111100011001010001000011"),
("101111010100010101010001110","101111011000010011010101001","101111011100011100001001111"),
("101111100000110111111111000","101111011011100101111000000","101111011001010011001111001"),
("001111011010111101110111110","001111010111001010111010001","001111100010100111111110011"),
("001111100011010000111011010","001111001000011111110100000","001111001111101011010110110"),
("101111100001001000100100100","001111100000001101011001011","001111010000110101100011110"),
("001111100010001110101001110","101111011100101101010111111","001111010101010111001000001"),
("101111011000000110100001001","101111001111101000101110010","001111010000001011011000101"),
("101111010010011100000110001","101111010001010011101011011","101111100010001001101000000"),
("001111001101110110011000001","101111010111111110011010011","001111011001010000100110100"),
("001111011001101111100001010","101111100000000111111111101","101111100000011100110110110"),
("001111011111111110110001011","001111010000101011111111101","101111011101011101110100101"),
("001110111110111000110101111","001111011001011010100101001","001111000011010010000001001"),
("101111100001010011100000011","001111011011010001101110101","101111011110010001010011000"),
("001111011100010111110010000","001111010011000100010101000","101111011010001001100101001"),
("001111011000010100101111111","001111011001101011100001111","001111011110110111000000110"),
("101111100010110010101110001","101111001110111001101010001","001111011011011101110000000"),
("001111100001010000101110011","001111010110101010011101001","101111010100011111001001010"),
("001111100001011101010110111","101111011011001001110100100","101111011100001110110010100"),
("101111100000111010110111111","101111100011010110001101101","101111011101010000100000000"),
("001111011100010010110010001","001111100011100101011111111","101111101000100011101110010"),
("001111000111010011010001000","101111011011010101101001110","001111011000111110010001000"),
("101111100011101011101011111","101111100000101100001010010","001111100000010100111011010"),
("101111100000001101010011110","101110111010111100011111010","001111010100011010101011011"),
("101111100011010100011011111","101111100011100000101110110","001111011111111101010101010"),
("101111100011101000101001001","101111100010010000001011100","101111011101110011011111010"),
("001111011100100100000110001","001111011101000100100011001","001111100001010001001011001"),
("001111011011100000111001000","101111011111010101010110110","001111100010111001010101011"),
("101110111010001101110101110","001111011100101000100110101","101111011100011100010101110")),
(("101111100001110011000101010","101111010101111111111001000","001111010110011010100101110"),
("001111010011101111100101101","101111100001111011011011001","101111011000000011110011111"),
("101111011111100011000111111","101111100000010111011100000","001111000001011011000011100"),
("101111100010100100111100010","001111011101000100100010011","001111100100000000010100011"),
("001111100001100101001011011","001111001110010011111111110","001111011011010010100100001"),
("001111011000100001000101000","101111100000101001110100111","001111100101001000100111001"),
("101111011001010001110011011","001111011101001101110111001","001111011000001001100100011"),
("101110101011111011110010000","001111011111001001100010000","001111010001110011001100111"),
("001111010110100100011110000","101111001111010101110001011","001111011000010100100111010"),
("001111100000111111000001111","001111100010010010100001101","001111011110111101100001000"),
("001111011110001110000001000","001111100110100110101011100","101111011010101000010101010"),
("101110111111101101000101000","001111001011100101110011110","001111010010010011010101100"),
("101111011000100010011111100","101111010001100000100001101","001111011101110000110010100"),
("001111100000010101101011110","101111010010001010101010101","001111011000010010100101101"),
("001111100001000011011111011","101111100010000011010111001","001111100001110100011101000"),
("101111100000100110111110010","001111100011110001000000011","001111001101010000001111101"),
("001111010101110111010010110","001110100101110100100101110","101111010001000000110100101"),
("101111011100101001000000011","001111100011011100010010001","001111011110000111001011100"),
("001111011011111001110001010","101111011011110000010100101","001111010100101000111101100"),
("001111001110000000100011000","001111010100010111100000000","101111010110101111100100111"),
("001111011001111110010111011","001111011011100100100000100","001110111101111110010001011"),
("101111011011100110101011110","101111100010101001110110011","101111011101011001100100011"),
("001111001000000101111111001","001111011011101110110011010","101111010011001100100001101"),
("101111100001101111110101011","101111001000001110110000000","101111100010001011001111000"),
("001111011100100010101110001","001111011101001001100001001","001111010001011000010110101"),
("001111100001001000010000010","001111100000001101110001010","001111100011111101011100010"),
("101111001111110001010001000","101111100000110111110011101","101111100011100110110100100"),
("101111100001000111101011011","001111011010110101101011101","101111000100111111000010010"),
("101111010001011011001110111","001111011100010101111011000","001111100100110010101111001"),
("101111100010011101001011010","101110110001100100010100110","001111100100111001011001010"),
("101111010011000111001101101","001111101000001011100101000","001111010011101110000101101"),
("101111001111010000000111001","001111100111011001110111010","001111100011100001000111110")),
(("101111011111001100001011100","001111100011010000101111011","101111011101101001011111010"),
("001111010000110110011011110","101111100010100010101100001","001111100000100010101001011"),
("001111001001001110011100001","101111011101111110011011010","101111100000100101011110000"),
("101111001001100000101000010","001111011011111111111000111","101111000101111000011100100"),
("001111010101101010011011100","001111011111110010001000011","001111011111110011111100011"),
("101111010010000101000111100","101111010100010001000010000","101111100000001001011000001"),
("001111100100110011110100111","101111011000011001100000101","001111100100111101011001100"),
("101111100001010001111100000","101111000000000010100111111","001111011000111000101001011"),
("101110110110010100111110111","001111011100111001101101100","101111010011000000010000000"),
("001111001100100111111110010","001111100011101111111111100","001111100100000011100010011"),
("001111100110100001010001101","101111000100011000100000001","001111100111000101111110001"),
("001111100011110111110110100","001111011010000111101010101","001111001010110001111010010"),
("001111100000011110010001110","001111100100010010100101001","001111011110001100011100111"),
("101111010001101001111010011","001111001110101100110100011","001111100011000001000010001"),
("101111011001110111001000100","001111011111010001011110011","101111001100111011011001111"),
("101111011100001010010111100","101111001101000010100000100","001111011000110100010001111"),
("001110111001000010010000001","001111100011000101011111111","001111010011000110101001011"),
("001111100100010000101101110","101111011001110111001001101","101111010000111011010100010"),
("101111100100010111110000010","101111100001010000100000101","101111011100010101111101010"),
("101111100010110111101010010","101111100011000010110011001","001111011000010110111001111"),
("001110111110010011011101011","001111001111000110000001010","001111100000011101110011000"),
("101111100010111010011111011","101111100010001101010000101","101111100000110011110101010"),
("001111011001001110000101011","001111001001100000111001010","001111010000111010100111101"),
("001111011110101101011111000","101111100011011010111010101","101111001100010111101010010"),
("001111100000110110100000100","101111011000111111100111100","001110111000010000011001000"),
("101111010010000010000110101","001111100010001101000110000","001111101000011000001110010"),
("101111011101010110011101111","101111010000001000001000111","001111011010010110110011111"),
("001111100101000111010010001","001111100010010101000010000","001111000010011011011111100"),
("001111100100101111011110111","001111100101001011000110110","101111011011011110100101010"),
("101111011011110010011100010","101111011010100000100110010","101111010000110100111001000"),
("001111010001110101100001111","101111011100101101101110110","001111010001100000101010010"),
("101111100000000001011010000","101111000110000101010110011","101111011010100001110101111")),
(("001111100011101010111101011","001111010101011000000111111","101111001101010111100111010"),
("001111010111000000011111010","001111000110101100001010001","101111100000101010100001111"),
("001111100011101110111100110","001111011000000010101010101","101111010001111010100011001"),
("001111100000000100110010110","101110110111100101011010001","001111100011000101010000111"),
("001111100101000001101101000","001111100000111011011010110","001111010111100100111000011"),
("101111011110100111001011101","001111100010001000001000111","101111010001001100110100110"),
("101111001010011011101000101","101111000001111111111010111","101111100001101111111111010"),
("101111011100110000100100010","101111100000001001110001010","001111011000011100110110001"),
("101111011100101101101001000","101111011000010011100101101","001111100000100111010111100"),
("001111001110101001111101011","101111010011000000001111110","101111001110111010000100110"),
("101111101000100000000000100","101111100001110100101000101","101111101000100110001101110"),
("101111001000100010100110101","101111010001011001101111110","001111010110100011000100010"),
("001111011101011111101101010","101111011001111011101001110","101111011111110101101111101"),
("001111011011110010000000010","101111011101010010001000101","001111010001101111110011101"),
("001111011001100110011001111","001111100010010101001100100","101111100001011010001011000"),
("101111001011001010101000100","101111011001100011000111111","001111011101101111010101000"),
("001111010101110100011011110","001111100000010011101011100","001111011000111010110001000"),
("101111100100111100000111010","101111010000001001110101011","101111011100110001000110110"),
("001111001010000001000110111","001111011101100110000101101","101111100011001111101101100"),
("001111001101100100101000100","001111011000101011010001110","001111011010010011110011000"),
("101111011101111011000011110","001111100101010011101101101","001111011010000110010011110"),
("001111010110001000100100011","101111100000010101011010110","001111011001011000101010001"),
("101111100011001010111010111","001111011000101000110100110","101111100001011110010100011"),
("101111011001010010100110010","001111100000101010100101110","101111100011000001001110000"),
("001111011010010010101000001","001111011000000101010110101","101111011010111001100111111"),
("101111100000111001100100100","101111011111000101100011100","101111100101100000100100010"),
("001111011011001101110100010","001111010111110001010001101","001111011000011110111100100"),
("101111010000110000000001001","101111100010111000010010101","001111010010010000001001101"),
("001111100010110100010000010","001111010011111001011001010","001111011011011110111101100"),
("001111001101011000100000001","001111100011101100000100001","101111010110011101111101100"),
("101111100010101101110100011","101111011001100010100010010","001111011001101100110001000"),
("001111000111000001011011001","001111011010111011000001010","001111100011000001100010010")),
(("001111010011101101000100001","001111100010011101011011010","001111010000001011111000101"),
("101111010111000110101110101","001111001001011001011111011","101111100001111011100100110"),
("101111011101000110111010011","101111011011100100101010110","001111011001011101011010011"),
("101111011000011010100011111","101111010010100101101011100","101111011111111010001011011"),
("101111100100100010101010001","101111101000000010011101010","101111010111000011001011100"),
("001111100011001001101010101","001111100011000101000101001","101111011101110101110001011"),
("001111011100011001110101010","001111010000110101101011101","001111011010100100101011010"),
("001111001001010011010011101","101111010010110111001110101","101111100000110001111101000"),
("101111100010010101001000011","101111010001011110101111001","001111100001100000000001101"),
("101111100001110101101101000","001111010011110100111110000","001111011101000100010110101"),
("001111011001101111010000101","001111011010111101000001011","101111011100100000100101000"),
("001111100011100111110101100","001111100001001110110100110","101111011011001100100101100"),
("101111011100001110000111110","101111100101001111001010101","001111100010011110011111111"),
("001111010001001110110110011","101111100010110010111100101","101111100000000100001010001"),
("001111011100111000011100111","101111010010100101100011010","001111011110001100111011001"),
("101111011111101000000101001","101111100000101111010010100","101111011101101100001101100"),
("101111011001001110101100011","101111011101011000110010111","101111011111011000001010110"),
("101111100000001001110101000","001111100001011000000101000","101111010110110011000100010"),
("001111000011111101011011111","001111100011010001101111111","001111100001111011111110000"),
("101111100000111110100101001","101111010100100101111110011","001111100010001110100001000"),
("001111010010100000000011110","001111100000000010101101110","101111000001111110101101001"),
("101111100010010111010111000","101111100000110101000110110","001111011110001111000101111"),
("001111011100111110001011001","101111000100011010010011010","101111001011110100111101100"),
("001111100000010100111001110","001111011010100001011010101","101111100001000110100001100"),
("001111011010011100100111010","001111011011110111110011110","001111100000000010101011011"),
("101111010101101100000101000","101111001001010000101011111","101111100000111101100001000"),
("001111010011000111010110101","101111011100100111000001111","001111100010110000011011010"),
("101111000101000010100100110","001111011110001001001110010","001111011010010101011010100"),
("101111011110100111011011101","101110101001010111011100100","101111011100101011110101000"),
("001111100000000000010110010","001111100010001011001011101","101111011011000100001111010"),
("101111100010010000111011010","101111011101111110110111101","101111100101111000100100000"),
("001111010010000000010110011","101111001110111111010011100","101111011101001000010011011")),
(("001111011111110001111110010","001111001100110100101110001","001111100100000000000111000"),
("001111011111011011110011111","001111011101111001101011001","101111011010100000110010000"),
("101111011111001010000111110","101111011011110000001111000","001111011101000000101011100"),
("001111100100110100100010100","001111011110000101011110100","101111011110111101011010101"),
("101111011010111000001000011","001111100011110011111110110","101111100001011101111000101"),
("101111011000001111001110111","101111001011110100111111110","101111011111100000000110010"),
("001111010111110100111101011","001111011110000001000010000","001111011001110000100011111"),
("001111011011101101100011101","101111100001001011011001111","001111100011110010010000011"),
("101110110110100011011000110","101111010110000011001001010","001111011111101001100000010"),
("101111100000011000111001011","101111100001000101100001110","001111010001101111000101011"),
("001111010010011001000111011","101111100001111100000010111","101111011100011011101001111"),
("101111000110001001100100011","101111100001001111010100011","001111011011100100001011011"),
("001111010010110110101101110","101111100000110001001101001","001111010111010101010101011"),
("001111100000101001100001010","001111100100101011101111001","001111100101001110010101100"),
("001111011110001101110101101","101111100000101111100000010","101111011110110110010010110"),
("101111011101010100100110111","001111100001101011101111011","001111100011001010111101001"),
("001111100010000011110010010","001111100001100110011001011","101111011011011101000100100"),
("001111100010010000001111010","001111011110011110101011011","101111011110000011111000111"),
("001111011000101101111010110","001111001101000010111110101","101111100000010001101111110"),
("001111100010010011111101010","101110111001011110011101010","101111010110110110110100111"),
("001111001000001101100010001","001111100000111100111001101","001111010110101001010000101"),
("101111100000110100111100001","001111001110110011100100000","101111010010111100101111101"),
("001111100001010101011000010","101111001101010110010001101","101110110011001110110100011"),
("101111100000001111111000110","101111100010101111000010000","101111000010110101000011110"),
("101111100001111010110010111","101111001010000011011011000","101111100010010011010110010"),
("101111011101110100101110011","101111001000111010001110000","101111100101100011101110000"),
("001111001000111010001011101","101111011111111111010000001","101111001011010000101111111"),
("101111011001100011110000110","101111011001010110011111001","101111100101010011111100110"),
("101111100100010001010001101","101111001111111011011100110","101111011111101001010100010"),
("001111011111000111111100100","101111010011101110000101110","101111000110110011100101100"),
("001111010101100111010111110","001110110011111001010000001","101111010011100101111101101"),
("001111011100101001110110010","101111001100111001111101100","001111011100000000110000001")),
(("101111011101100000101001001","001110110001100000100111010","101111011011110110111010000"),
("101111100000001001010010110","101111011100110110010111111","001110110001000100010000000"),
("001111001110000000001101011","001110111101100111001111001","101111010001001110001001000"),
("001111100001101011001000010","001111100000100110101001110","101111010101000110110101010"),
("101111010101110001111101000","001111011011001100110001101","101111010000011111010001011"),
("101111100100000010100111011","101110101110000011010100100","101111011010010111000000010"),
("101111011101010001011110000","101111001001001001000110101","001111100001100001100110110"),
("001111011011000101111101011","101111100011010011111000111","001111011110111101001111111"),
("001111100010111010111011100","001110101010001100010101011","001111100000110101100100000"),
("001111101000110011001000111","001111100100100110100001100","101111010001110010011111100"),
("001111100010100101101101101","101111000000101111111110011","001111101000011100011110100"),
("001110100011000100011000001","001111010100101110110001011","001111011110111100101000010"),
("001111100000010110001110001","001111100101001001010011010","101111010101010101111111110"),
("101111100010100100100010110","001111000000110011010010011","101111000010010101011011000"),
("001111011011100110001000101","001111011110111000110010110","101111100010100010010001101"),
("101111100001001010100011000","101111100010100101100100010","101111100110111100100101110"),
("101111011110101100000001000","001111001001010100100100000","101111010000010111000101010"),
("101111011111001101100001011","001111001100000001011101100","001111011100101011100101110"),
("001111000100110101101110011","101111011100111001111111110","101111100000100100011000010"),
("101111100011011101100110010","101111100101001000111010010","101111011010101101101101110"),
("001111011010100001011000010","101111100000110011001101001","001111011100100010111110001"),
("001111000011111110001001010","101111100000001001000101001","101111011011010010010111001"),
("001111100011000111001000001","001111100000001111000101101","001111010101100100011110010"),
("101111100001010010000011110","101111100011011111111111110","101111011000111110010110011"),
("001111001101010010001111011","101111011000110100101100010","101111100001110111001000000"),
("001111100101001010110011000","001111100011001110000101011","101111011001110001100010010"),
("001111010010001100110101000","101111010011011100001111011","101110111011001000010000101"),
("001111011000010101010010101","001111011101001010110101111","001111100001111011111100111"),
("101111001011100001000011101","001111100000100000111100101","001111011101111101010111010"),
("001111001001111110111111010","101111100001001010100011100","001111100000111110111000111"),
("001111011001110011011110010","001111001100001111010001100","001111100011100110100101101"),
("101111011011101101111010110","001111100011100101111001001","001110111001010011110010100")),
(("101111011100011110010111011","001111100010100110100000110","001111010001001000111000101"),
("001111000000010100100110001","001111011011101000000111000","101110111111011101111101101"),
("001111001101110101100010011","101111100011110011100010101","001111100101001001110100011"),
("101111010100011011011111110","001111011000100000001110100","001111100000011011111001101"),
("101111100001001011100111001","101110111110100100011100111","101111100001110010101101001"),
("101111011110010110100011010","001111000001011110001111010","001111100000101111011101101"),
("101111100110011101010011010","101111100101001101010000000","001111011101010111111101010"),
("001111000001110000011111000","101111010100000111011000011","001111011101111011110111010"),
("101111100010111000101010110","001111011011010111100100011","001111011111100100001100110"),
("101111011010101100101100000","001110110011000001101011100","001111011100101100001000010"),
("101111100010001010010100100","101111001010000111101110111","001111100110000000000111011"),
("101111010001110000011011010","101111100110011100101110110","101111011111001101011010011"),
("001111010011001111110000101","101111011110110110111011000","101111010000000100100101101"),
("101111100110100110101100100","101111100100100100011110010","101111010011001111010101001"),
("101111100000001000100101101","001111100011001101111000011","001111011011110001110110110"),
("001111000000010110011101111","101111011110110111100111101","101111100100100011010110111"),
("101111100001110011110110010","001111100010011110111110111","001111011111011011100110100"),
("001111011111111010010010100","101111000000010010010111010","101111011111100010101000010"),
("101111100011100011001110001","001111011011010011000111010","001111011110011111101011110"),
("101111100111101101110101010","101111010001110001100000100","001111100000010010000001101"),
("101111010110001010000011101","001111010100000101110001010","101111100101011100000011111"),
("001111011110100010101000011","001111011001001010001100011","001111010110010100101010011"),
("101111010111101001110001010","101111011101100011101010001","101111010110001011100001000"),
("001111010000100100000101101","101111011110100111001010111","001111011001011010000100110"),
("001111001110000100000111000","101111011110110001110001111","001111011001110110110100111"),
("101111001100110000100010111","101111011110011011110001101","101111001100001000100000101"),
("001110101010000011110011101","101111100010000011001011100","001111001010100010101101100"),
("101111011110100111110101010","101111011011111010110001101","101111011000100000101101001"),
("001111011110010100001011000","101111011111110110111101100","001111011010110001000100010"),
("001111100100011001101011011","001111010001011001010011010","001111100001011100111001010"),
("001111100000001110111001000","001111100000011101100111111","001111010111111101110100000"),
("001111011000011111000111011","001111011010010001011110001","101111100001000011001110110")),
(("101111011110000000011001011","101111001111001001110111011","101111011001100000100010110"),
("101111001000001011100111100","101111011110000000100100010","001111001101100010110000010"),
("101111001000111000000010001","001111100001101000001111011","101111011110111111000000010"),
("101111100001111011100101001","101111100011010010011000001","101111010101111000111010110"),
("101111011111001000100110111","001111100001010100001111010","101111100010010110100010011"),
("101111100011010111001010100","101111011001011110000001101","001111001101100100101011001"),
("001111011001010100010001100","001111010000010111011100011","001111001110011111000100011"),
("001111001001111111001011110","101111010101000111101001000","001111100001011000110100111"),
("101111011001000111010100010","101111011010111011110000000","001111011101111111100011001"),
("101111000100001100100000000","001111000011011010101011101","101111100011100110101110001"),
("001111100011001001000011110","001111100010101110110011100","101111001101110110011011010"),
("101111100000100101000100100","001111011101001011101110101","001111100000001001100111111"),
("001111011101111110010110101","001111010011100001000100000","101110110010011101111100101"),
("001110110110011100011111101","101110011110011110110001110","001111001111000001001010010"),
("101111011011011011110001101","001111011100000100011100001","101111011011100101101100111"),
("001111100000111010011011100","101111000101011011101100011","101111100001110101011101110"),
("101111100010000001011001010","101111001011011101010100101","101111010100001000011000101"),
("001111001011101010111011100","101110001100000101110010011","101111011101100011111111100"),
("101111010111000010010110001","101111001100110011110110101","001111001100100101011011011"),
("101111001000100110101100000","001110111011000111100100111","101111100000111000000001111"),
("101111100001001101000111110","101111010111111110001100001","001111011001101011110001001"),
("101111011110100111010001001","001111011010100000010111100","001111001110101000111000111"),
("001111011001011011111101110","101111011111101001110000110","101111000110110110111001001"),
("101111011010111010100110000","101111011010000101101110101","001111011001000000111010011"),
("101111010110000000000100111","101110111111000110011010111","001111010101110000000011011"),
("001111100010101000101000110","001111001010010111011010001","001111001000111000000111101"),
("001111011011110100100000001","001110111101101111101100101","001111000111001111101110001"),
("101111011011000000010010010","101111011011100110011011110","101111100001010101110011111"),
("101111011010001011011100010","101111010011111001000011001","101111011111011011011011011"),
("101110011100100011101001101","101111100010111011001110010","001111011000000111110001010"),
("001111100011001010001010110","101111010000010100001000000","101111000110001111011010001"),
("101111100010010110101101000","101111100010101111111011000","001111011110110110011111010")),
(("001111011000000110111001100","101111100010010111110001100","101111010100000011110011101"),
("001111100000100011011110100","101111100011011110000100110","101111010100111010011101010"),
("001111011011110010111101110","101111010001101000011101001","101111011110000011101000110"),
("001111100001000101011101110","101111011101110010001001010","001111010101011010110000111"),
("101111100010011011101100001","001111011010001010011001111","001111011001001011111100101"),
("101111100000011000000101001","101111011010110101111010010","001111011111010101000000111"),
("001111010111001101000011000","101111010010011000001011100","001111100011110001101101101"),
("101111100000010010111011011","001111011101111100111000000","101111011010101010101000000"),
("001111011101111000000101110","001111010110100000101001110","101111001001000010011110011"),
("001111011111010011111110111","101111100001001000011000000","001111010011011000101100001"),
("001111001110011101000011110","101111100010100010111011011","001111100000101000110011111"),
("001111100010101000101100110","001111011111000110000010001","001111100100100111011001001"),
("001111100010101001110010101","101111011100001010100110110","101111010101001111001000101"),
("001111011100011110011110011","001111010000100100110111000","101111001110100110100101100"),
("101111011110001000101001101","101111011011100111001000100","001111011010100000110000011"),
("001111010011010011100100111","001111011001111011001001100","001111100010001011100110011"),
("001111100010000100100110001","001111011101111001001110010","001111011111110000010111111"),
("101111100011101101011011000","101111011101101100011010011","001111100001000011011000110"),
("001111010010011000110001101","001111010101100001110001100","101111001001101011011101101"),
("101110110100010111111011000","101111011000011000011010001","101111010111111111000000110"),
("001111100000010111101001011","001111100000000111011001011","001111100000101010010110110"),
("001111100000110110101000011","101111100001111000011110100","001111010101000100111110010"),
("001111000111110110001001010","101111001011010111110001001","101111011010010010000101000"),
("101111011101010101101000010","101111100100110000011001101","101111100000110101011010110"),
("101111000011000100101100110","101111011111011010101110010","101111010110010001100001100"),
("001111100000110110101010101","001111100010001101110101011","101111001101100010111001010"),
("001111100001111000001000100","001111011010100100100010100","001111011011110000010101000"),
("001111011100000101001100001","001111010000000011111011110","001111100010111101110110011"),
("001111100000111011100100000","101111010001111011011011001","001111010100011111100101010"),
("101111001011100111100101010","101111010101011111001100010","101111011111011111000001001"),
("101111011011110100001001100","101111011000010111010101100","001111100000000010001001010"),
("001111100000000000000011000","101111011110010111101011110","001111001111111100111000100")),
(("101111010011111111101001100","001111000000011101110100000","001111100100111100001111011"),
("101111010010100001101101110","001111100001111110100111000","101111001001001110111000010"),
("101111000011101010111100101","001111100010000000010001011","001111100001010011010010100"),
("101111001111001011110000101","001111100011100111010111000","101111010011111110101100101"),
("001111011110001010000111001","001110111100100000111110000","001111100000101100101001001"),
("001111010001001000101111100","001111000001110101000001101","101111011110101000011110111"),
("001111011101101111000100111","101111000111011010101011000","101111001100000111010011101"),
("001111100010010001110010100","001111100010100110011010110","101111000000011011111100010"),
("101111011000101000011101010","101111010111011000011110110","001111100001101111110010010"),
("001111011111000101101001001","101111001110110101000110101","001110101001010101010000110"),
("101111100001101011011000001","001111001010010101001101000","101111011110001010101010110"),
("001111011111111001010100111","001111011110011001101000000","101111011111000001101000100"),
("101111100001001011110011011","001111000010000001011101010","001111011001100110010101111"),
("101111100000101011100111111","001111011000011111001111001","001111011011101110011101010"),
("101111100010000100001001110","101111010000000111101011001","101111011101101101011110111"),
("101111000110111110111000000","101111011001000111001010101","001111100000001011001100110"),
("101111010101111011000010001","101110111000001000001100011","101111011101100101000011110"),
("001111011111000010010100011","101111100000000110000001011","001111000110100001111110101"),
("101111100100001110101001101","001111001010100101010001011","101111000100111110000010101"),
("101111100010110000101111000","101111011011100010010001000","101111100001001110000010011"),
("001111100001001011001011001","101111100000100101100110010","101111010010111001101000001"),
("001111011111010011001111111","001111100001100101011111011","101111011010010000001101111"),
("101111100101000111111000010","001111001011001101100101110","101111000000101101100010010"),
("101111011110111000010101100","101111011010111011101101010","001111100001011011101000000"),
("101111001111000010111100111","001111010010010001110001101","101111100000111110011000101"),
("101111011000101100110001111","101111000101000100010101101","001111001011001110110011000"),
("001111100000001110011111110","001111010110011000101110100","001111010010001000000100011"),
("101111011110110000001100100","101111011010011110001000001","001111100011001100110101010"),
("001111100011010001011111111","001111011101100110101100011","001111011111111000111011111"),
("001111011111011101010100111","101111010000101010100011010","101111011011110011111010111"),
("001111011011111101010110101","101111010100000100001010111","001111100011100000010010110"),
("001111100110111000111100010","001111101000101011110000101","001111100001001111001010000")),
(("001111001001011110110111100","101111100000011101011101000","001111000001111001100011001"),
("101111001001001101000001011","001111100010101110001010111","001111010011011001101010000"),
("001111010000111011000011001","101111011111101110011011001","101111100010011100100000100"),
("101111011101110000110010111","001111100000111111000000011","001111100001010011110110100"),
("101111100010011011101110000","101111010011000001011001101","001111100001010001000011001"),
("101111011110110100001011001","101111100010010110111010001","101111010000010001101111001"),
("001111011000000000001011001","101111100100011000110001001","101111010001110111110011010"),
("001111010000110111001111101","101111100010000101101111110","001111010000110111100011010"),
("101111011110101101110101001","101111010011010101010111010","101111011111110101011101000"),
("101111010110010010100010000","101111100000010001100011101","101111011100000011001001110"),
("101111100011100110100100111","101111010000100101000000011","101111011110110110110110110"),
("001111010100001110111001110","101111100001000111000111100","101111100000110011100100100"),
("001111011111101010001000011","101111100010000011101110101","101111100001010010101111000"),
("001111011111100110110000100","101111010011100111010011100","101111010100101110111011100"),
("001111011010100010100111001","101111100010011110100111110","001111011100010100011100010"),
("101111011011110000010000011","001111011101110010010010111","101111100000101100100100001"),
("101111011110011101001001000","101111001001000110101101111","001111011101100010110101101"),
("101111000010100000010000110","101111100010101111100100100","001111001001100101101010111"),
("101111011101110101001100011","101111100010110011001000001","101111010001001001001101100"),
("101111011101011110110110111","001111100000010011101111110","101111011000011001100100001"),
("001111100011001001000000101","101111100000010111111011001","101111100010100110010011001"),
("001111100010000011001100001","101111001111000101110111111","101111010101111010101101100"),
("101111001001001010000010111","101111100010111000001110010","101111001001000001110010010"),
("001111010000011110110010001","101111000011110101011111001","001111010110100110001111100"),
("001110111100010101000110011","001111011100100011111110101","101111010001001110011010001"),
("001111011110110110011111100","001111100010110010011100100","101111100000101010011010100"),
("001111100000001011111010111","101111100010001010000101000","101111011100000000000000011"),
("001111100000101000001001101","101111011111110111010011100","101111011001111100101111110"),
("101111001011110101100010011","101111100001011110000100011","101111100010000110010011000"),
("101111011000000101010001000","001111011111000000111110110","101111100001101010111011001"),
("001111100001110101011010101","001111011001000010111101000","101111011111001001101000111"),
("101111010100111100111010100","001111100010100000010010000","101111011100011000010000111")),
(("101111001000000000001100110","101111001001000011011001110","001111011001101100111001010"),
("101111011110011001110111001","001111011101100010011111100","001111010001011011101000000"),
("001111001001011110100110011","101111010111001001010010000","101111011010101001000010101"),
("001111011110111101100100110","101111100000010111011011001","001111001011001001000101110"),
("101111010011110011101011011","101111100010111001001011010","001111011011101100010111000"),
("101111001001111000100100100","001111100000000101010000010","101111011001101111110000101"),
("101111100010010110100101110","001111011100111110010100100","001111011111000010101010101"),
("001111100000011100011001000","001111010100000101010011000","101111011101001110011100010"),
("101111011001000110100010011","101111010000100101011110110","101111010001010101001111011"),
("101110111100100111011100110","101111010010110100101100011","001111100010010001110010000"),
("101110111001110011100111110","101111100010001100111100000","101111010101001111111000101"),
("001111011111100001100110100","101111010101011110011101011","101111100000100110001011010"),
("101111100010101110010011010","101111011011010000101011010","001111100001010001000101011"),
("001111011010111100110100110","101111011000111110011111101","001111011001001000011011111"),
("001111010001110001011001110","001111010011100010011101001","101111100100000011100110110"),
("001111011000000001110011111","101111011001001110110110100","101111010000010110010010110"),
("101111100011101100011100010","001111011010111011111000000","101111011011100011000011101"),
("101111011000011000011110001","101111100011110111000110111","001111011001011100010001111"),
("101111011011010011001100010","001111011100101100101100110","001111100000011111010111001"),
("001111010001100101111001000","001111011101011001100001111","101111100011000000110011010"),
("101111011010101010000100101","001111010011001000001001110","101111011001101110000011111"),
("001111011110111001101001111","001111010000110100011000100","101111010001101001010011111"),
("101111000100100010111111110","101111100010001011010110110","101111100010100100000110111"),
("001111011100110100001101111","001111100011100000000101101","101111010111101010000000011"),
("001111011010000000010001110","101111100000011000111100011","001111011000011110011111111"),
("001111100011011000100101000","101111100001000001101111001","001111011101100011110100010"),
("101110110010011110011111101","101111001110011111000111110","001111011010010010111011100"),
("101111010001010011101001110","101111011001101111010011010","001111010010010100110110000"),
("101111001110011001111101010","101111010111000011111100001","101111100011000011110110111"),
("001111011110011111011100101","101111000110001010001011001","101111100001001111010111110"),
("101111010111111101011000111","101111011000101110110000000","001111011100011010111110101"),
("001111010001111100010000101","001111000101010011000111001","101111001010101010100010111")),
(("101111100000110001010111100","101111011111111110001011000","001111011111111111001011001"),
("001111011111111011010101000","001111010011111000101100001","001111000010011001101100010"),
("101111100010000110110011110","001111011011011110110100111","101111010111001101101000011"),
("101111011011111101011000101","001111011010000100010111101","001111001110110000100010010"),
("001111100001011010001010011","001110110100000001110001000","001111100101101000101101110"),
("001111100001100011100001101","001111100101011010011010100","101111010011110100100110000"),
("001111011110100010000111100","101111010010111111000001110","101111001010010001011000111"),
("101111010001110010101110000","101111010011110011110001101","001110110101011100011011001"),
("101111100010101110110010110","001111011100010000011001100","001111100101001011000001001"),
("001111100000101000101000001","001111100001011111010010000","001111010001011100011101111"),
("001111011110110011010000001","101111011101011100001000001","001111100000111010100001100"),
("001111100011010000111010100","101111011010000010111001001","101111001100100100010000100"),
("101111011001001011110000001","101111000010010100011100100","001111011101011000010110001"),
("001111100100010111010010001","001111011111010100100010101","101111100001100001000100111"),
("001111010100010000011011110","001111011100100111011000111","001111001010101111111111001"),
("101111010011111001110010001","101111100010000001111001000","101111010000111011000001011"),
("101111000100000010110001110","101111000101000111111111111","101111100001101110101000000"),
("101111010110110000111010011","101111010011000111110101111","101111001000000010111111001"),
("101111100101011001110110010","101111100101010010001111001","001111010011001010010100110"),
("001111100000001011101101001","101111001010011111111101011","101111011000101011101101011"),
("001111100010110110010111000","001111100011011000110000001","101111011010101001011111101"),
("001111100001000000111011001","001111011011011010000000110","001110101001010000111111011"),
("101111010110010001001010001","001111100110001101110000101","001111100011110100001010000"),
("101110110000101100101101100","101111100010111111111000101","101111100010011010110101011"),
("101111011100011110010010010","101111100000011011010111100","101110111100011110001100001"),
("001111011111101000001011101","001111000110110011001001110","101111010000111000100101101"),
("101111011001011101100100010","101111100001000001000110111","001111100001000011101100000"),
("101111011100001010110000111","001111011110110111100010001","001111011100000000111100001"),
("001111100111111001011000101","001111100000110010011101101","101111010010110011001100101"),
("001111100000101111100110001","001111011111111110011111111","101111011011101000011110011"),
("001111101000001000100001010","001111100011101000101100010","001111100111011111001010100"),
("001111100001010110100010111","101111000000100010101110011","101111011011111000001100111")),
(("101111011000000111110111101","001111100000100001010111001","101111100000010110010011010"),
("001111011011001011010111000","101111100011011101011001101","001110110010000010010110011"),
("101111001011110100100000111","101111001100011110010110111","001111010100100111101000000"),
("101111000010001000111111011","001111010011110000011011010","101111010010110011100101100"),
("101111011110001001100011010","101111011010101100010111001","001111010111110110010111101"),
("001111011011000100001110110","101111000010010100011000100","101111011110010101010011100"),
("101111101001001110100000111","101111100111000101010100011","101111011101110110010101011"),
("101111001000110111101010111","101111010111111111011010000","101111011011110011010101100"),
("101111011001110100100000110","101111010101011101000011001","101111011010111001010100011"),
("101111010001111100001111001","101111011111110110111111000","101111100100010001000100100"),
("101111010110111110110000100","001111100000000001010100110","101111011000110011111110100"),
("101111010011100000101111110","101111010011100101000010001","001111010110000001111110011"),
("101111010000101110110001010","101111100010000100111000001","101111011101011001011111011"),
("101111010110000001101001111","001111100001000001001110101","101111100011100110000110110"),
("101111011011011101111100100","101110100111010100100111000","001111100000100000110000010"),
("101111010010110011001001000","101111100110010011101101110","101111100101001110001100111"),
("101111011100000111010011000","101111011010110011111101010","101111001010001100110011100"),
("001111100100010001000101111","001111011001100010010111111","101111100010100000101111001"),
("001111100101000101101011101","001111100001100000101100010","101111011011110001000111100"),
("001111100100000101010001111","101111010010110000001110111","001111010011101101001001011"),
("001111000101001001001100100","101111011000000011100100110","101111010010101110010101011"),
("001111011011010100110111110","101111011101101111100110101","101111100011100101011011000"),
("001111100010000010010100101","101111100001100100001011000","101111100000110011001000110"),
("101111011110000000001111111","001111010010010111110000010","001111010100100111101001100"),
("101111010100100101011001000","101111100000101110010010001","101111011010000100111100100"),
("001111001010100110000101101","101111011111110000010001101","001111001111100100111101101"),
("101111100011101111110001000","001111010000010001110101100","001111001101110010100111001"),
("101110100000101011101000101","001111010100001101000110111","101111011100110100000010000"),
("101111011111011101110010011","101111100100111110000000011","001111100000001001101001000"),
("101111010101111000001110111","101111101000001000100000000","101111100000001000110000111"),
("101111100100001000101110000","001111011011101100110100101","001111011101110111011000000"),
("001111010000001011100001010","001111000110011111000101111","001111011100110001101100110")),
(("101111001010000001001111110","101111100000010101101001111","101111011011110000100100110"),
("101111011110011011010000111","001111011101101100100111001","101111011110001110111001100"),
("001111011111000111100001110","001111011100100011100001001","001111010110110101111100111"),
("001111010010001100110010100","101111011010010011101000110","001111000001100000111010010"),
("101111011100110011011010100","001111100100011100010111110","001111010000110101110001101"),
("101111011100001111101110010","101111100000000111111111110","101111100001001001101000111"),
("101111010100001000011010111","101111001010001101001110000","001111100101000110101101111"),
("101111011011111010111000011","101111011100010011011110000","001111000111010101101010110"),
("001111011100010010111110010","101111011111101111110011110","001111010110111110010101101"),
("001111100101001100100100101","001111100011100000110110011","001111100100000110110101001"),
("001111100010010111100100110","001111100011111001010100101","001111011011100100011011001"),
("001111100000110000001010110","001111001011000001001011000","101111000000000011101011111"),
("101111011000101110100011001","001111011001000100001010101","101111011101001110111101101"),
("001111011101010001111101111","101111000110000110101111000","101111001101101010000100100"),
("001111100000101100010111000","001110111110100001110001011","001111100000100101111111101"),
("101111011011000000001110000","101111100000011101000110101","101111001000011010111011001"),
("101111000001100011110010001","101110100000110110011100111","001111011010001010010101100"),
("101111100001111101101101001","001111011100010001010010010","001111100001011011001101100"),
("101111100110111001111010000","101110101000111101111111010","101111011110000111010101101"),
("101111101000000010010101101","101111011000010010100101011","101111010111011011111010001"),
("001111100001110100110000000","001111011010100001110101010","001111010000111101110110010"),
("001111011100000001010110000","101111010111110101100011100","101111000101000011101011001"),
("101111010111101111010111101","001111010110001011001001100","001111100010001010101111101"),
("101111100011101110010010100","101111011000011100011000001","101110111100101001100101100"),
("101111011100110011010110010","001111001110110111011001111","101111011001101010101110010"),
("001111100010111110110011011","001111100011100111100100001","001111011101110010110001110"),
("101111010111101001011101101","101111100011101101000011011","101111010000000010100110110"),
("001111011110101001110111111","001111100011110001111000000","001111011100000000011001100"),
("001111010100001001111101000","001111011100001110011011000","001111010011001010110001110"),
("101111100010011001001000100","001111011000001100010101111","001111011101000111100101001"),
("001111011011110011000001111","001111100110101010110000010","001111100111001000110001011"),
("001111000001110111011001000","001111011100010101100011101","001111011000010111000001110")),
(("001111100011111011101101110","101111100010100101100101010","001111100010001001100011000"),
("001111011011100000010110111","101111001100111011100000011","101111010111111111010101001"),
("101111100010011101001001100","001111011111111000100100110","101110110010011100001000010"),
("001111011110110001010000010","001111010100101001111000101","001111100001111110010110000"),
("001111010100011000011001010","101111100000010000000000111","101111100000111101100111111"),
("001111100001000001010111010","101111010111010001101010000","101111100000111010011111000"),
("101111011001100111010000110","101110111001000000110001000","101111011001010010111111101"),
("001111100000100011011011101","101111100001000000111011111","001111000101111010101100110"),
("101110111001100100010011111","001111010101110010010001011","001111100001100111000011001"),
("001111100000000110010000011","101111011100011110010001011","101111011001100101000011001"),
("001111100001100001001110101","101111010011001011100011100","001111100100000010001100110"),
("101111100100000100110000000","001111010111001010011011100","101111100100101001111010001"),
("001111010110010101110001101","101111100010100000101011011","101111010110100111010001011"),
("101111011001100010110000110","101111100011000110101101000","001111010110011111011001110"),
("001111011011110111111001010","001111010001100001000101100","101111011111101010111111100"),
("001111001010111110011111101","101111100001100001000011000","101111011110000000001010101"),
("101111100001110010011100001","001110111011000001011110001","101111100000011000100111110"),
("001111100000001010000110000","001111011001100100011011011","001111100011011101101110111"),
("001111100100110111000000011","101111010100000011011101011","001111100101011010101011111"),
("001111010101001011110010011","001111100001011110010111010","001111011010101101111110100"),
("001111011000111000011010101","101111100110100010001100110","101111011110010011001011110"),
("001111011100011111010000000","101111100010001111011011000","001111011100111101000100110"),
("001111001110000111111000100","001111100011101110101100011","001111100101110111010110011"),
("101111100000000101011110100","101111100001101101110100100","001111010001111000101011001"),
("001111011000010010100011010","101111010110100101110111110","101111011110010110000100010"),
("101111011100011110110011100","101111010011001100111011111","101111011101010101011111010"),
("001111011010000101101101101","001111010010101010000101000","101111010111111101011000000"),
("001111011101010011110010010","101111011000010010010111111","001111100001110000110001000"),
("101111010100000011010011001","101111011101011100110011010","101111100010101100010010101"),
("001111011011111110101010101","001111001111101011001110100","101111001111010011101011100"),
("101111100001110010100010110","001111011101001010011101001","101111010000110101011000101"),
("101111011010101111101010111","001111000100100001110000110","101111100001101101011011001")),
(("101111011111010111010100101","001111010011010111001001001","001111100001110001011110001"),
("001111010111011001010110010","101111001100010011111001110","001111010011001010011111010"),
("001111011100110110011111101","001111100011110111100111011","001111100010010101010000001"),
("101111100000001111000000000","101111001000111100100000101","001111100000010010111111011"),
("101111001101011010100111000","001110111000100000110000000","001111100000011100001010010"),
("101111011101001000111010011","101111011111000110101000011","001111100010101000101001101"),
("101111001001010001100111000","101110110001011100011011010","001111100000011011010110011"),
("101111100001010001000110010","001111011111110001110110100","101111100011001010111011001"),
("101111010011011010110110110","101111100010111010111111010","001111001010001000100011111"),
("001111100000000010111110001","001111010000010110101011001","101111010110000100010000110"),
("001111100101110000110000111","101111011100111010111011000","001111011100100101011111000"),
("001111010100110110001011101","001111001100010100001001111","001111010010011001100010001"),
("001111010010100111100011011","101111100010000000111111110","101111100011100100000100101"),
("101111010011100000010110100","001111011010010011101101111","101111010010100011011111110"),
("101111010100001100000001011","101111100000001001011000010","101111010100101000010101000"),
("101111100010100001101000011","001111010111011001100100011","001111100000011100011010011"),
("101111011110000100001000100","001111011011001100010011111","001111100000001101100101100"),
("001111100011010110100010011","001111001001000000010001100","001111010000000011001001010"),
("001111011100001111111100101","001111100010000011001010100","001111001000011101110001001"),
("001111100000110000010111010","101111001001001110111110110","101111011000011101101101110"),
("001111010001011010100001101","001111011010010101011011111","101111011111110000101000100"),
("101111100001001100101101010","001111100000011100000011000","001111100010001100101011011"),
("001111011011111111101101001","001111011011010010010001100","001111011011001101001110111"),
("101111010100110010100100101","101111100001111110000001010","001111010000100100010000101"),
("101111010011101010100100101","101111100001110000001110101","001111011101010001001001001"),
("001111100001110011010110000","101111011000010001101000010","001111100011011000111000000"),
("101111001010011001101100100","101111100000101000000111110","001111011000000110000101011"),
("001111100011111111010110001","001111001010111101100011001","001111100000101000111111111"),
("101111000101100011110101000","001111011101101010011101001","101111010101001110101001010"),
("101111100000111000010001100","001111011010101101101010110","001111011111111101010011010"),
("001111001011011100001000010","001111101000010010101000001","101111010110011101110101101"),
("001111000100101011000001011","101111000110000010011100011","101111010001100111001100011")),
(("101111011010010010001110111","101111100010101010110000100","001111100001111000010001011"),
("001111100001000011010111010","001111011010011000000011001","001111001100110100010000000"),
("001111011111011010010010101","101111011011000101100001010","001111011110011011011101010"),
("101111010010000100010100110","001111100001001111100110010","001111100100011001100001010"),
("001111011011000111011010000","001111001101101110001011000","101111011000001000011110001"),
("001111001111111001011110001","001111100100110100101101101","101111000010110011101001101"),
("001111100010010010101000110","101111011100101111100011100","001111001100011110101100010"),
("101111011011011110110111011","101110101011101100101111111","001111100010101010000010101"),
("001110111011001011001101101","101111100000101111110111010","101111010010111001100110111"),
("001111001011111011111111000","101111011001111100000100001","101111011011110100000011010"),
("001111010010110101010111110","101111100010100101011110100","101111100011001011110111010"),
("001111001111011010001010101","001111010111111010110101111","101111100011011110011110100"),
("001111010001001001101110100","001111010010111111110100101","001111011001101111110001001"),
("001110100010001110111000000","001111011101001100100011001","001111100011100001111111000"),
("101111010111011101000100000","001111010110001000100010011","001111100000101011101000011"),
("001111100000000100011110100","001111001011100010110011110","001111011010100101111000011"),
("001111001110011100001000111","001111100000101110000000010","101111100001110111010000101"),
("001111000100000001000001001","001111011010110000010111011","101111010000100111110101010"),
("001111010101001100110100011","101111010110100001000110111","001111011011111110100100101"),
("101111100010000111010100101","101111100011011110111110000","101111101000000011111101011"),
("001111100001100001000011000","001111011010011100110100010","101111011110101010010010001"),
("101111010101101010011010110","101111011101010010011110000","001111010000000100101000100"),
("001111000111111011100010111","101110101101111000100110101","101111100000001001110011010"),
("101111001010010011000101110","001111011010111010010111001","101111011001101001111001010"),
("101111001011010110011110101","101111011100110011110111000","001111011001011010100001001"),
("101111011000000111001000100","101111010001001100111101110","101111100011011101010010010"),
("101111100110101110111010010","101111001011111010011101101","101111000101110010110010010"),
("101111011100101000000110100","101111010000110111011101011","101111010110111101110000110"),
("001111100000101000011110011","101111011000001110011111011","001111011010110011100010001"),
("001111011111011110100100100","101111100001000100000001011","101111010000001000011010101"),
("101111001010111100110110101","001111100000001010111111101","101111010101111000100001011"),
("001111101000101111010000000","001111100111001101001100001","101111011000101011101001011")),
(("101111000100010011111011010","001111100001101111110100111","001111100001101110111100011"),
("101111010111000011000000001","001110111111000000001000110","001111100100111011111100111"),
("001111001001101101100010011","101111011011101000111101010","001111100101010111101110010"),
("101111001000000011100001111","001110111101100011111010100","101111011000110100000001100"),
("001111010001110111000000100","101111011011010010110001010","001111010111100000101010100"),
("001111100001100100110000000","001111010111101101000010101","001111000111001111010111111"),
("001111001011011101101011100","101111010011101001000110110","001111011111100011011100101"),
("001111001101011000110100001","101111011100111001100001001","001111010110000010111110110"),
("001111001001101111110101100","101111010011011010000001000","001111100011000100001100100"),
("101111011111001100101011110","101111100101111111100010011","101111100100100110101111010"),
("001111011001100011110011110","101111100011100100110000111","101111100100011111101110000"),
("001111001010100111111111111","001111011010111110101001101","001111011011101001101010111"),
("001111011010100100011001100","101111011101111110000111100","001111100000111000111111011"),
("101111100010000101011111011","001111011111011001010010001","001111001010110001001100011"),
("101111100000110011100110101","101111011111000100110110111","101111100001011011111010101"),
("101111011111100001100111101","101111100000011011001111011","001111010011111011111010100"),
("001111010000010111000001011","001111010100101101000110001","001111100000101000111101100"),
("001111011010011101101011110","001111010001111110111010001","101111100011110110000000111"),
("101111100011010011101101011","101111100001001110001101010","101111100010000100001000000"),
("001111100000000000010011000","001111010011001011010000111","001111100010111111100100110"),
("001111100000110101000001001","001111011000110000101010101","001111100011001010110101000"),
("101111011001010011001110011","001111011000011010100110111","001111011101100111001010001"),
("101111011100111111100001110","001111000011110111101101011","101111011100100000001000000"),
("001111010100101011100101100","001111010101010100111110001","001111100100010000010100110"),
("101111100010010001000000110","101111010001001000010111110","001111100001100101011001101"),
("101111100001000110110110100","001111010000110101111000100","001111100000010111111000100"),
("001111011101000000111000110","001111011100100011100100000","001111100100011111110100100"),
("101111011011110100011010000","101111011101110110011111001","001111100000101111111110101"),
("001111010001101101001000101","001111100000101000111001001","001111010110110100111011111"),
("001111010010100000110110000","101111011111110101001100100","001111011010100000101010010"),
("101111100010011000101011011","001111001000001101011010000","101111100011011110011111101"),
("001110100110100001111111011","001111001111110110011011001","001111001111001111110100110")),
(("101111101000000101101110000","101111100100110001110000100","001111011011000001001100011"),
("101111100000010001111110110","101110100000111100101100101","001111011001110010100100010"),
("001111010001100101100111111","001111010011010111110010000","001111011010110111101001001"),
("001111100011111101001010010","101111011001011010010000001","001111100000100110101011100"),
("001111100000111101000101101","101111100010001111101110001","001111001100110101110010001"),
("001111100100111111010000100","001111101000000101100100010","001111011111001010001110110"),
("101111100011011011010001111","001111011110100000101110101","001111011111100000001110101"),
("101111011101101111000100100","001111010010001011010000010","101111011110100010101100110"),
("101111100001000111010001000","001111001100110011001011101","101111011111110011101000000"),
("101111010001010101111001000","001111011010000100111111111","101111010011010000101010001"),
("101111100000101010110100100","001111011011110001101001010","101111011100110100101010011"),
("001111010000011110000110101","101111010001011110111001011","101111011010111001011100111"),
("001111000101101101111111101","001111010100101111000001100","101111011111011010100100100"),
("101111100110110010101100011","101111100001000111111011001","001111100001101010000001000"),
("101111011111000111001101001","001111011100100101000101101","101111100001101001101111000"),
("001111010011100011010110010","101111010101010100001001000","101111011111000001100101011"),
("001111000000111101110111010","101111011110010110101101000","001111100001000010110110001"),
("001111100001000101111101101","001111100001011101000111111","001110111101001100010111110"),
("101111001001011111001111100","101111010110000000001001110","101111100011101000101001101"),
("001111001010011000001011011","101111100010101110010010000","101111100010011011010110011"),
("101110010011000000001011000","101111011110111101110110100","001111100010010001110001011"),
("101111010111000110001101111","101111100101000100010101001","101111100001101101011000000"),
("101111011110110001010101100","001111001110100110111000001","101111010100011111011100010"),
("101111011000001100000011011","101111100101011010101101101","001111011001111011111101000"),
("001111010000001001101111100","001111010010111011110001111","101111100001110100010101011"),
("101111011110011101001001100","101111100000010101100001011","001111100011111001110101010"),
("101111100101110100110011110","101111100000100000001011010","101111101000001000101110101"),
("101111100000000111111111101","001111011101000000111100110","001111011110011111101101001"),
("101110101101010000101000000","001111001110110100100000110","001111011111011101101001010"),
("101111101001011011101010101","001111001111111111000011011","101111011100101001110011010"),
("101111011010010100001110111","101111010001010011000100001","001111010000001110111001000"),
("001111010001011111010010111","001111100110000001111110010","001111100001001000001101010")),
(("001111010000100000111000011","101111011000011101110110011","101111011001011011111100011"),
("101111011110011000100100010","001111100010101010001010100","101111100001001111100110000"),
("101111100010100011000010101","101111011101110110011110110","101111011001110010000001101"),
("001111100100000010001010010","001111011110101010001100110","101111100010010001001101011"),
("001111011010001100000010100","001110111110100001010111101","001111010100010000011011101"),
("001111100101000011100110010","001111011001111001010110011","101111100010011111011011010"),
("001111011000001001011010001","001111100011110101001101110","001111010101100011010001110"),
("001111001101001001111000000","001111011111000010100110011","101111010000100001100101010"),
("101110100111001010111001100","101111011011100011000000010","101111100001010001100110100"),
("001111010010001010010001000","001111011010110001010111111","001111100010010000001010101"),
("001111011101110000011101100","001111011010101101011100100","101111011000111101110100000"),
("001111010100011111010110110","001111011100010111100011010","001111010001001111010001010"),
("001110111101001101100010100","001111010011100100010000101","101111011001001010111001011"),
("101111010011100011011100101","001111100001001100011010000","001111100010000000001001101"),
("101111100010011000100100111","101111011111000100111011011","101111101000000010110011101"),
("001111100101100111011100001","001111100101011110011110101","001111011011111001011011000"),
("001111000011111111011101100","101111000111110000000010010","001111011111001010011011010"),
("101111001011001001110100001","101111011100101110100100000","101111010001111100001110100"),
("001111010101100110001100000","101111100001011000100011001","001111100010110101111011010"),
("001111010111110110110011100","001111100000111010100110000","001111100011010111000101010"),
("101111011111110110111010001","101111010111000011010100001","001111100001100010000101111"),
("101111010001001001110100000","101111011000000000111000001","001111000111011010111010000"),
("101111100000101111010110011","101111100010101001011000011","001111011100010000000010111"),
("001111100101110111111000000","101111010000011111110100011","001111100011001101111100001"),
("101111100001110100110111111","001111011011110000001000111","101111011011111001001001111"),
("001111100000000111111001011","001111010000110111101010001","101111100001001101001000011"),
("001111000000000101010000100","101111011100101111100000110","101111010101010011100000101"),
("001111010010010111111110011","001111011100110010100101000","001111011010010010111111001"),
("001111100000000011110111011","101111011001110100010001101","101111100010001101001100110"),
("001111100101110010011101101","001111011011111000111110101","101111011111101110110100010"),
("001111011000011001011000100","001111100100011001111101000","101111010110001110011111000"),
("001111100000010101010011011","101111010000110001001100111","101111100000110111001111101")),
(("001111010000101001001111101","101111011001000010011000101","101111010111101001111100010"),
("001111100001101011111000110","101111010011010010101001101","001111011010000100101001010"),
("101111000011101100000001110","001111100000011100111101110","001111001101100000111101010"),
("001111010110011110100011111","001111100010011010100010111","001111100101010011000110011"),
("001111100000001011011101110","101111011001110011110101001","001111100010000100001101101"),
("001111100100100011101100010","001111001011111000110110111","101111011101110010010000011"),
("101111011111010001110100001","001111011010011001111111000","101111010011001110111101001"),
("101111100001101000001101101","001111010001001111101111000","101111011011111001100100100"),
("101111011111100011011111111","101111001010101011010000100","001111011100110111011010100"),
("001111100101011110011010110","101111010001011001010110111","101111100000100000111001100"),
("001111010000010111000110100","001111100110010101110001101","101111010011100110011001110"),
("101111100001100101101110001","001111011011101111111100000","101111010110011111111000110"),
("101111010100010110001110000","101111010010110011000100010","001111000011000011110100000"),
("001111011001110110001100110","001111010011101010110110111","001111100000001100010110100"),
("101111011111101010100101101","101111010101110100110111111","101111011011111001100100101"),
("101111100011111100100101001","101111010101110111000011101","101111001111010011001010110"),
("001111011101000010110110110","101111100010000101010100101","101111011011100111101111110"),
("101111011101111000110110000","001111001000011100100110111","001111011011000101010100010"),
("101111100001111111100001011","101111100111110101010000101","101111001100110001100011100"),
("001111011100000111101111100","101111011000100110100000111","101111100001000010101101010"),
("001111011101011010011111110","001111100010110000001011010","101111100011001010110100001"),
("001111000101011100000000110","001111001000100000000001010","001111100001010101110010100"),
("101111010111111101111011101","001111001010110100111110110","101111010111100101111000101"),
("001111000111000001100011111","101111001100001000010010001","101111100010111001011111001"),
("001111010100001001000111001","001111000011011011010001010","001111011110011000010100111"),
("001111011000000001111100100","001111011101111101011000011","101111011000001101001100011"),
("101111011101011100111110001","001111011001010101100000001","001111011000100101100011111"),
("001111011001011110011011111","001111100001011011010101111","101111011101100111000010011"),
("101111100000000011111010101","101111001111100001110110011","101111100001110110010110100"),
("101111011011001010011100101","101111011011101010000011101","001111011100111101010110000"),
("101111010100101100001010000","001111100100101001000010000","001111011010010100100011001"),
("001111010000001000110000011","001111011010101011111111001","001111011101000100011101100")),
(("001111100000000100100100111","101111010010101111110100001","001111011110011111101100000"),
("001111100011011111011101110","001111100011001110100101101","001111011000010101110111011"),
("001111010111110010011010000","001111010011001101010001011","001111100010101111010110010"),
("001111010010010001010100110","001111011001011100110101100","001111011010100101000000010"),
("101111011000000100001000010","001111100000010111101101101","001111100000100001101100000"),
("001111001110100111011000011","001111100100000000101001110","001111011110100101011111001"),
("101111011110010010110001011","001111010000000101010100010","001111100101001111001101100"),
("101111100000000010101110000","001111011011011000000010011","001111100010110111110100010"),
("101111011100100110111110011","101111100000110000001000001","001111100000010110101111001"),
("101111001001111101111110001","001111010011100010100110101","001111100001111101100110010"),
("001111010001101010001111001","001111100100100111010111010","001111100100110101000010101"),
("101111100000011001001100101","101111011101001011010010000","101111011111101000001110000"),
("001111011001110111100111101","001111010001101110100001101","001111100110110010101010000"),
("101111010011110010111011111","001111100000111101001010010","001111100000100101011000110"),
("001111011000100110000110001","001111100011010000110101101","101111010111110101111011110"),
("001111000001110100001000111","101111000010001110111010111","001111010100010011001101000"),
("101111011010000000000000101","101111011011111010101101110","001111010010111010111110100"),
("101111011010111000101110001","101111010100001001001111000","001111001011111110101100000"),
("101111100100011000101001110","101111100011100111110010100","101111011001000010011100101"),
("101111001101101000111000101","101111011100110101111111110","101111100000001110111100101"),
("001111001001000001010111000","001111010110010011010100100","001111011001001111111110100"),
("101111011000000100110101101","101111011101011100011011000","001111100100000100010100000"),
("001111100011000000011110111","001111011011000100000000111","001111010111110001000000001"),
("001111011110110011100001110","101110111101011010101010000","101111100011101000110000101"),
("001111011110000011110000000","001111010100100001011011001","001111100010111110010110011"),
("101111001101110101100100110","101111010001011001101101111","001111100011100101100110010"),
("101111100011011010110110100","101111010111111011111111001","101111100000011111101110100"),
("101111010100001000011100100","101111011010001000111011000","101111100000000101001100110"),
("101111100000110110001000101","001111100100111101101111011","101111011111000100100010111"),
("001111011000101110010010101","001111010001000110011110010","001111011111100010010000000"),
("001111010111100100000111111","001111010101011111100110010","101111001010110100011010000"),
("001111011011000101110010100","001111100010101011110111100","001111101000010011111100101")),
(("101110101101110101001111001","101111100000010101111000010","001111100100000101000111000"),
("001111000010010100111011010","101111011011010110000110010","101111010100110011111001001"),
("101111010101111001100111101","001111100011011101011100110","001111100110110101001110100"),
("101111100001100111010000101","101111100011011110010011110","001111010000001011001100011"),
("001111010011111011011100011","101111011110101000110111000","101111011111111100100110000"),
("101111011101011100011110101","101111100101011100101000011","101111001001110011101101100"),
("101111011101111000010010011","001111010010000101000011011","101111011101100001110101101"),
("101111011001100110101001011","101111011000011010111100010","001111011101000000101010000"),
("101111100010011100010001011","101111001111010110100111000","001111100011010000010000011"),
("101111100000101111100111001","001111011110011001011101101","001111011011111110010110111"),
("001111100001011011010011100","001111000110011001000000001","001111001000000110101001100"),
("101111001110100110110100010","001111100001001010011110010","001111100101101111011001010"),
("001111010100110111100111111","001111010100010110111111101","001111000001101110111101001"),
("101111010011100110110010111","101111001001101011111000001","101111010100101011000010101"),
("101111100011101101111110110","101111011010110101000011100","001111010000000111011101110"),
("001111001010101110011011000","001111100010101010001110010","001111100000100011110000100"),
("101111011101010101001011000","101111000111101010100010001","101111100010011011000110110"),
("101111011000101000011111001","001111010100101111100110001","101111100001010000110101110"),
("001111001101110000101010101","101111100000001000101110111","001111001011110110011011011"),
("001111000000010110001010010","101111011011010101011100110","001111010101110001101010111"),
("001111001100001100101111100","001111100100011001010111111","101110111001111101100101000"),
("101111011101100110010111001","101111100010100001100000011","101111011001011010111100111"),
("101111100000110011001101001","101110101101001101101110000","101111001111110110000000000"),
("101111011001110110001111111","101111011110000001101011101","001111011100100011101111101"),
("001111010100001010011101010","001111010110000110001001010","101111011110000001011110100"),
("001111011010001101100110000","101111011000110010110110100","101111011001011111010100001"),
("101111010001001111110110000","001111100010110110010011000","001111100101111001111001011"),
("101111100010110101010110101","001111000011010101111001001","001111011101011111111000100"),
("101111100001011110000011010","101111001010001011010011101","101111011000000101110100000"),
("001111011101101000111101011","001111011100010011111101101","101111011001011010100000011"),
("101111100011010101000111001","001111100011000010001111110","001110111000110110001111110"),
("001111100100010010001010011","101111100010101010000101000","101111011010010011110011011")),
(("001110111011010111001101010","001111100000001100000010110","101111011101010010011010110"),
("101111011010101000011110010","101111100001110010000110101","101111001101001111001000001"),
("101111001010001011000001011","001111001110001001001100101","101111011101111010111101000"),
("001111010010101101110101000","001111100100000100111111011","001111100000111111100100101"),
("001111100100101010111000100","001111100011111000100110110","001111100101101100010010000"),
("101111010010010100111111101","001111100011111011101110100","001111011110001101001110101"),
("001111100100111000110111000","101111100000011000001000000","101111001010000100100110100"),
("001111100010111001100010001","101111011101011001100010111","101111100010000010011110010"),
("101111011000100100010100101","001110111010101100001001101","001111100001000000010100110"),
("101111010100110000110101000","001111100000001111000100100","001111010010011110110010111"),
("001111011010000000100001101","001111100011100000011110001","101110111000101111110101001"),
("101111100000101111101000100","101111010010001000111101101","101111011001100100011000101"),
("001111100010110001001010001","001111011001101110110101110","101111010100010100101100001"),
("101111100011001110101101000","001111011000100000011111110","101111011000111011100111000"),
("001111100001110111011011010","001111011001000001010110101","001111011110011111011001100"),
("101111100010100001101010010","101111100001111111010011110","101111011001101101010100101"),
("001111100010000100001000001","101111011000001011011110000","001111100001101001110101101"),
("001111100010110111101000100","001111100000001101000000001","101111100011001001011000101"),
("101111100010010011001010110","001111011000011001100100100","101111000101111110110000000"),
("101110110011110110011101000","101111010101010011101000100","001111001110111011100111111"),
("101111011010011100111010000","101110111110111000010100010","001111010010011100001001000"),
("001111001111100011111001000","101111011101110100111000001","101111011011001000111100000"),
("001111100001010101100101110","101111100011001000000000111","101111100001100010011010100"),
("001111001000011000101001011","001111011001001111000001100","001111011101101010000011011"),
("101111001000000000111101101","001111010010001111101011110","101111010001100111001001000"),
("001111100011001000100111011","001111001010000010111010101","101111010101011111000010110"),
("101111100100001010000101000","101111011010111110010001000","001111011111011001110010111"),
("001111100001000110010001110","001111010001000101001111000","001110101000000100000110000"),
("001111011000111010100111000","001111010010000010010011010","101111010001001000101000101"),
("001111001000000010110110111","001111100011000110000100011","001111100001011000101010101"),
("001111011000011110001001011","001111100010111001001010011","001111100011110000111101011"),
("001111100011001010001101101","001111011011000101111011100","001111011110010000101000101")),
(("101111100010110101101010000","101111011000111100101000011","001111010101110010001000010"),
("001111011010110100011010111","101111010110001100011001000","001111010010101010000100110"),
("001111011101010000000110100","001111011110001001111001011","001111010111111110011110010"),
("001111001010100101001110111","101111011000000000111101110","101111010000011011011111100"),
("001111010101100001110010111","101111011010100011110010111","101111010101001100000000111"),
("001111100001110001100110011","101111010110101011100100111","101111100001100010110101100"),
("101111011000000100110000100","101111011011011010010100100","101111100001010110001110010"),
("101111100001010111011001101","001111010100101110010100111","101111100010011011010010110"),
("101111010011101010010000000","001111010100100011100111101","001111100000011111110000011"),
("101111001101100010111110000","101111011011000000011000101","001111011101110101010001010"),
("101111001001011010100100101","101111011011111001110011011","101111011000010101100110011"),
("101111011110010010101001010","001111010101110110011101100","001111010111000001010101100"),
("101111000011111100000001010","001111010101011110101111111","101111001010010110000100001"),
("101111001001000100111000111","001111100000001000000100101","001111011100010101111001000"),
("001111100010000011011110001","001111001110010110100000011","101111010000001010001001111"),
("001111011011000000100001110","001111011100111100101011001","101111010110101001100100010"),
("001111001011101001010111111","001111010010100000101001101","101111011101011101001101011"),
("001111011010101000111111101","101111100001110001011110010","101111100010101001011011001"),
("101111001010001011001011111","101111011001011010100111101","001111011000001100001001101"),
("101111011100010001010011111","101111100010100100101011110","001111001111110001001111000"),
("101111100001100111111001110","101111100001010011010001000","101111100000011010111010001"),
("001111011111111111001100010","001111100001100111110100000","101111100000110000001000101"),
("101111100000000011001000000","001111011010110101111111110","101110110111010111111111001"),
("101111100010110001001001000","001111001110100011101000101","001111100001001100011101001"),
("001111100001000010010011001","001111001101010110010101101","001111011101001010001001011"),
("001111011111001001110011100","101111100010111011101110000","001111100001010100110011111"),
("001111011011001010000011001","101111100001100001000100111","101111010001011001010011111"),
("101111100000110100110111111","101111010011101111001011101","001111011010101101100010110"),
("101111011011110010110110101","001111011111010101100000110","001111011011011010111100001"),
("101111100011001000101000110","101111100010111110101010001","101111011000111101011111011"),
("001111011010010110001101001","101111010010110000010111100","001111011011001110010101001"),
("001111010100110011101110010","101111100000001110010110011","101111010000001101111100010")),
(("001110101011010000100101010","101111100011001010011101100","101111010010001100010110001"),
("101111100010100011101010001","101111100001100100010001000","101111011011001000001110001"),
("101111011111100011101001111","001111100100111101100110111","001111011000101111010001100"),
("001111100001110100001011101","001111001100010001010110110","101111010001100010001101110"),
("001111010000100100101111110","001111100011001110010110001","101111011000111001110000111"),
("001111010010000101111001011","101111010000101001011000111","001111100001001101110011111"),
("001111100011011100100011010","001111000011000010101001001","101111011110000011011111101"),
("001111011110101110111111101","101111100000101101001110010","001111100000101010000101101"),
("001111011101001001101101001","101111011011011011000110011","101111011010011011101000011"),
("101111011101100101010011100","001111010101101110001101001","001111100001010000010111011"),
("101111010110111010011010110","001111011010011101000111101","001111001111011010100000011"),
("001111011100011000001110111","001111100100000101100101011","101111011100110001010010110"),
("101111010000111101000101011","001111100101011011001100001","001111001000110011001010110"),
("001111100000010100111001100","101111010000000001000010010","001111100011100100001011101"),
("001111011001010100100011111","101111011110100011010010101","001111100011101001111011010"),
("101111100011010000110001010","101111011111101000100111110","101111011010011110000110011"),
("101111011011101111110010000","101111001001011001010110000","001111100010100100001000101"),
("101111010110000110111010001","001111011111101001100101001","101111100001001011101110111"),
("001111011011110100000100010","101111011111001111111010010","101111100001010011000100011"),
("001110111010111111100101100","001111011001010111110011100","101111011000111010100001100"),
("001111100011011011100100001","001111100010000101011100111","001111011010000101110100100"),
("101111100000101001001100001","001111000110000110001011110","001111011110100110011000110"),
("001111100011110101101111110","101111001001010010000101101","001111010101011011011100100"),
("001110101111101001000001110","101111001100111000100000001","001111011101011011110011111"),
("101111001011010000011110011","101111010011110101111110000","101111100010111111110111001"),
("101111011100010110101000110","101111010001101000101101010","001111100011101011101001111"),
("001111100011110010100111111","101111011111000110101101110","001110111100110111001110010"),
("001111011011001101000000011","101111011011001101010110100","101111011110001111000101100"),
("001111100110010000101001001","001111100001010010100110010","001110110001111011010010011"),
("001111011110101011011111100","001111011000111110001011101","101111100010011101110001010"),
("001111100001011000011110000","101111011011010100110110011","101111011000111000111110000"),
("101111011001011100110001100","001111000011000011000100100","101111011111001110111001010")));

end fpupack;

package body fpupack is
end fpupack;