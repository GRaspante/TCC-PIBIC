----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 05.08.2023 00:18:30
-- Design Name: 
-- Module Name: cnn_conv2_c_tb - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_unsigned.all;
use IEEE.NUMERIC_STD.ALL;
use work.fpupack.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity cnn_conv2_c_tb is
--  Port ( );
end cnn_conv2_c_tb;

architecture Behavioral of cnn_conv2_c_tb is

component cnn_conv2_c is
    Port (  reset_conv2 : in STD_LOGIC;
            clk : in STD_LOGIC;
            start_conv2 : in STD_LOGIC;
            samples_conv2 : in in_Conv2;
            filter_conv2 : in filter2;
            bias_conv2 : in biasConv;
            ready_conv2: out STD_LOGIC;
            output_conv2: out out_Conv2);
end component;

signal sreset_conv2, sclk, s_start_conv2, sready_conv2 : std_logic;
signal s_samples_conv2 : in_Conv2;
signal sfilter_conv2 : filter2;
signal sbias_conv2 : biasConv;
signal soutput_conv2tb: out_Conv2;

begin
uut: cnn_conv2_c port map (     reset_conv2       => sreset_conv2,
                                clk               => sclk,
                                start_conv2       => s_start_conv2,
                                ready_conv2       => sready_conv2,
                                samples_conv2     => s_samples_conv2,                                    
                                filter_conv2      => sfilter_conv2,                                
                                bias_conv2        => sbias_conv2,                                
                                output_conv2      => soutput_conv2tb);
                                
clk: process
        begin
            sclk <= '0';
            wait for 5ns;
            sclk <= '1';
            wait for 5ns;            
        end process;
        
stimulus: process
    begin
        sreset_conv2 <= '0';
        s_start_conv2 <= '0';            
        wait for 10ns;            
        sreset_conv2 <= '1';
        s_samples_conv2 <= ((others =>(others => (others => '0'))));
        sbias_conv2 <= (others => (others => '0'));
        sfilter_conv2 <= ((others =>(others =>(others => (others => '0')))));
        wait for 20ns;
        
        sreset_conv2 <= '0';
        wait for 10ns;
        
        s_start_conv2 <= '1'; 
        sbias_conv2 <= secondConvBias;
        sfilter_conv2 <= secondConvfilter;
        s_samples_conv2 <= (("000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","001111000111100111001010010","001111010000011011111110111","001111010111111100111010110","001111011001010010110001111","001111011011110001101101000","001111011100111101100000111","001111011110011111111101001","001111011100110011000001010","001111011011110111000111101","001111011001000111001101000","001111010110001100100010101","001111010100110101111111000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000"),
("000000000000000000000000000","000000000000000000000000000","001111010110001000001001101","001111010110000110111001111","001111010101000110101001011","001111010110001110100110110","001111010100111110011010000","001111010101001000011100110","001111010100110110000000000","001111010101100011111101010","001111010101111111001110001","001111010100001001000011110","001111010011110110010010001","001111010100101110011011101","001111010100100010001100011","001111010011100101101011111","001111010001100111110110111","001111010001010101100111110","001111010011001110000000110","001111010010110100011011111","001111010100111010010010110","001111010100101000100010001","001111010011011001011100101","001111010010110111110000110","001111010110010000010000101","001111010100010001011111111","001111010101111000010001100","001111010110001011110100100","001111010101011010101100111","001111010110010101011011000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000"),
("000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","001110001000100001010000100","001111010000011000011011011","001111010101011100101100110","001111011000111100000100000","001111011010111010110100111","001111011100110110100110111","001111011101000011100010110","001111011100011001110111001","001111011011110011011100110","001111011001011111101110110","001111010101001100010000000","001111010101100011011110111","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000"),
("000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","001111000000011011010010111","001111010010001110110111100","001111010101100000010010011","001111011010001111101100100","001111011100100001100110000","001111011111111110100010001","001111011111001000111110010","001111011110111101111101001","001111011100001101100000000","001111011010001000000101111","001111010110001010111011111","001111010001001001011001100","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000"),
("000000000000000000000000000","000000000000000000000000000","001111000111101101011000110","001111001110101000011000001","001111001101011110001010001","001111001011011010110110111","001111001100001101000101110","001111001110001001101011001","001111001011100100000010000","001111000111101111101011100","001111001011111011100101111","001111001110101101001110100","001111010000000111111100100","001111010001001110001111111","001111010100000100100010011","001111011000011011000011101","001111011000000000000010100","001111010110111010110011110","001111011000010000111111010","001111010110110110001010000","001111010100001000111100100","001111010110100110011000010","001111010110000000011100110","001111010101111000111111101","001111010011011011110111111","001111010000111000010111000","001111010001111000000111000","001111001111100111100011100","001111001011101011111101100","001111001111101001110000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000"),
("000000000000000000000000000","000000000000000000000000000","001111011000000010010010010","001111010111011111001111111","001111010110001001101000000","001111010110101101101000110","001111010110001001111101000","001111010110101101101000110","001111011000000010011000000","001111010101111111000110110","001111010101001000100010000","001111010100110011011000010","001111010100000001110110011","001111010100110000000101100","001111010011011101111110000","001111010010011010100000000","001111010100101100101011011","001111010011111101101001000","001111010100110000111110001","001111010111001001110111100","001111010111101010010010101","001111010101110011001110101","001111011000000100011010100","001111010111011111111010111","001111011001010001011110100","001111011001000110010111101","001111011000101101011100101","001111011000101111111111110","001111011001011011110011101","001111010111011011010011001","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000"),
("000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","001110110100011101001011100","001111010001011000000101001","001111010100000101111000011","001111011000110101111111100","001111011001100000011100011","001111011011111111111001101","001111011011100111111010000","001111011011010000101000000","001111011000110011010101101","001111010111010010100101010","001111010010100110101111010","001111010010011001010101100","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000"),
("000000000000000000000000000","000000000000000000000000000","001111010001010001101001000","001111010010011001010001011","001111010000001110101010011","001111010010000100110101110","001111010001001010110011110","001111010001010110010010110","001111010011100010000010001","001111010101101001000101100","001111010011101011101010101","001111010001000000101001101","001111010000010100100001110","001111001101011101101000100","001111000110011001110000111","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","001110110101000111111010001","001110101011000110011010010","001111001000100000000000111","001111000001001000111010001","001111001010000000010100011","001111001000110000111111001","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000"),
("000000000000000000000000000","000000000000000000000000000","001111000110100100111001111","001111001111100000001101110","001111010001100000010001011","001111010100010001011110110","001111010101010010111001110","001111010111001111101001101","001111011000111010111000100","001111011010010110010100101","001111011011010001100110011","001111011010111111010111010","001111011010100000111001100","001111011001110011111010001","001111010111111110001111110","001111010010111011000011100","001111001001110100001010011","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000"),
("000000000000000000000000000","000000000000000000000000000","001111011001011010101001001","001111010110011101111001001","001111010100110111100101110","001111010100110110101110001","001111010011011110000000001","001111010011000100110011011","001111010010011110100101001","001111010100001000100000001","001111010001111011010001011","001111001101100111011001100","001111001101010000010111010","001111001101101111011101011","001111001110111011001001111","001111001011000000000101100","001111001010111110010100010","001111010001011010111111110","001111010010101011100101101","001111010100000110100100011","001111011000110010111001011","001111010111111100001011101","001111010111111010110110101","001111011000001110010001110","001111011010101111111000111","001111011010011111010000101","001111011010010111110111110","001111011010001111100110110","001111011010011100010010111","001111011001101110000101011","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000"),
("000000000000000000000000000","000000000000000000000000000","001111010100011100001101101","001111010110011111001101000","001111010011010001110000111","001111010100001011000100110","001111010100111110000110000","001111010011111001000000010","001111010100010100011011100","001111010100010100100010111","001111010100110110001011101","001111010011000000001101111","001111010011101110001101001","001111010010001101011000001","001111010010000000100011001","001111010010011001111011010","001111010001100101101001010","001111010001000100000100110","001111010001111101010001011","001111001110001000100011111","001111010010110100010010100","001111010010000011011001100","001111010010100111010100000","001111010010010110101101110","001111010001011101001101010","001111010100000011110110011","001111010101101101101010000","001111010011111111000001000","001111010011101100011100000","001111010110010010000111001","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000"),
("000000000000000000000000000","000000000000000000000000000","001111010100111010001011011","001111010100100010101101111","001111010011001010010001101","001111010100101001000001101","001111010100111100010000101","001111010100010011110101110","001111010100001100011001110","001111010110101011100110110","001111010111110001010011011","001111010101001011011001100","001111010101111100101001100","001111010101000111110011111","001111010100101010011100110","001111010010111000101110101","001111010000100000110000000","001111010001000011101101110","001111001111010110110011111","001111001110000101010000000","001111001110110000111001011","001111001100001111110011111","001111001101000100110000110","001111001101011111101110110","001111001000101001100101010","001111001111100001011001010","001111001111000000101010001","001111001111111001011110101","001111001101001001100101001","001111010010110111100111011","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000"),
("000000000000000000000000000","000000000000000000000000000","001111010110110000111000011","001111010011110101101111100","001111010100000100101000101","001111010011111000010001000","001111010100001001000000101","001111010011001100000001111","001111010100100001010001101","001111010100111000000100001","001111010011011111110010011","001111010001101010100111000","001111010001001111001010101","001111010001101000101100011","001111010000110101001011101","001111001101100011010111100","001111001101011010110000000","001111010001101100010111010","001111001110100001011111110","001111010011001101101000101","001111010011000111000101001","001111010100010000011010101","001111010001100110000111110","001111010110001000000100011","001111011000000011101000010","001111010101101011000010010","001111010110010110101000100","001111010100101110101000001","001111011000000010000100000","001111010101001000111010001","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000"),
("000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","001110101100011001001111110","001111001000111101011110010","001111010010100100101000000","001111010011101101011101000","001111011000011001010101100","001111011001011111111010010","001111011001010111000111110","001111011001001001010010110","001111011000110011010111010","001111010101001110110001100","001111010000110101011011011","001111010000110101000111011","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000"),
("000000000000000000000000000","000000000000000000000000000","001111011001001001110011010","001111011001100100111011110","001111011001101100101100010","001111011011010100110011111","001111011011100011011011010","001111011100000110111110101","001111011101011100110100001","001111011110101001000100010","001111011111011010111010100","001111011111001100000001011","001111011110111001000111110","001111011101111111011001001","001111011100111011001111101","001111011010010010011111110","001111011000001000001010101","001111010010100010110111111","001111010000001100100100010","001111000110100011101110011","001111001000011111000100000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","001110110011011011000111101","000000000000000000000000000","001111000000110110011011010","001111001001001111001110111","001111001110111100000010100","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000"),
("000000000000000000000000000","000000000000000000000000000","001111011000100010011101101","001111011000011011100100110","001111011000010110110010100","001111011000110111010011011","001111011000110100100101111","001111011000011110101000010","001111011001100111010001101","001111011001011101100110100","001111011001011010110101010","001111011001000000111010011","001111011001000000010101001","001111011000100011010001100","001111011000000001000100101","001111010101010000111110000","001111010100101000000000100","001111010010001100111101111","001111010011011101101111011","001111010010111101010001001","001111010011010000111110100","001111010010000001000110110","001111010010010000000011000","001111010001001010111101001","001111010011111011011111101","001111010011101000011100001","001111010100100011010101110","001111010110010110101101110","001111010101001111000110100","001111010110001010001101110","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000"),
("000000000000000000000000000","000000000000000000000000000","001111010000011011010011111","001111001111111101011100011","001111010000011011111101111","001111010000110110101111010","001111010000011110101111001","001111010000000101100101100","001111010000111010011111011","001111001111101011111100100","001111001110100101101000000","001111001111110101110011110","001111010000011010001100101","001111010000101111000010011","001111010000011001101001000","001111010001100111000010011","001111010001110001110110100","001111010010111000001000111","001111010010010010000011000","001111010011010100110101000","001111010001111100010000011","001111010011000100001100101","001111010010101101110001001","001111010101000101010000010","001111010001011011111101101","001111010010010101110111010","001111010000111000110111100","001111010010101110001001010","001111010000100100111101100","001111010010001011110111101","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000"),
("000000000000000000000000000","000000000000000000000000000","001111001010111110000111101","001111010011110100111101010","001111010110111011001000110","001111011000100110110000111","001111011010000101100111101","001111011011001010110000101","001111011100110110011111100","001111011111001110000011011","001111100000010111011011011","001111100000110001110110100","001111100000100111100001001","001111100000010000010011010","001111011111001001010101011","001111011011111001100110000","001111010110100100111001111","001111001011001100100100100","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000"),
("000000000000000000000000000","000000000000000000000000000","001111001001100001010100100","001111001001101101110011100","001111001000111101010111111","001111001010000010101111101","001111001011101001100110100","001111001101000100000110111","001111001100010011110101110","001111001110000011011000100","001111001111000100001000100","001111001111110110101000001","001111010000010101000101100","001111010001000100011011111","001111010001001000011011110","001111010000001011000101111","001111001010000011101000010","001111001100011000010111001","001111000111101100100010010","001111000011100001101011000","001110110100011010000010001","001111000000000001001001011","000000000000000000000000000","001111000000010101011001011","000000000000000000000000000","000000000000000000000000000","001110111001110110010100110","000000000000000000000000000","001110111001111001010101110","001110111100101011110111000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000"),
("000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","001110111101001010101010010","001111000000010001000100100","001111000101001111010100001","001111001010111011101100011","001111010000111101101011111","001111001011001111100001010","001111010000000000101001111","001111001001010010100110111","001111000011101001111011100","001110111101011001101111000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000"),
("000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","001110111001111011011011111","001111001011000101100011101","001111010000001001111000010","001111010011000011111011111","001111011000010000111100110","001111011001000111100100101","001111011001110110010010101","001111011000110100100010110","001111010111011001011000100","001111010100101001000111111","001111010011011100001100110","001111001001000101011011110","001111001101001010011001100","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000"),
("000000000000000000000000000","000000000000000000000000000","001111000101111000010001100","001111000011100111111101101","001110111011110010001100000","001110101101100001000100110","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","001111001001001001011111111","001111010000001000001001001","001111010011000111110110100","001111010110110111000100110","001111011000101010111001101","001111011000110001110101110","001111011010010110011010011","001111011010100001001011010","001111011100010110001111111","001111011011011000001100011","001111011010000001101111001","001111011010000110000010011","001111011000001101101000111","001111010110110110100010001","001111010100100111111001010","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000"),
("000000000000000000000000000","000000000000000000000000000","001111010000111101001001010","001111010011110010110100111","001111010010110000001100011","001111010010001001010111010","001111010010101101101110000","001111010011000000111010111","001111010001010001000101011","001111001101001101110001100","001111010000010001010111011","001111010010011111110000101","001111010010110100101001100","001111010100010100110111111","001111010111010010101100101","001111011001111101011111100","001111011010010100011001011","001111011010001010100011010","001111011010010111101011001","001111011010101100110101111","001111011001010101011110011","001111011010100010000011111","001111011010011000110011100","001111011011000101011011010","001111011000110111001101101","001111011000000011110100010","001111011000100011010100001","001111010110100010011000011","001111010110010010000000111","001111010101010101001011100","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000"),
("000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","001111010000101011111010001","001111010000011110110011010","001111010101011000111100101","001111010110011001100100010","001111011001111100101010100","001111011010000010100101001","001111011001001011011101101","001111010110001010011001010","001111010101111100000010110","001111010011001011010110111","001111001111101111010000010","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000"),
("000000000000000000000000000","000000000000000000000000000","001111010110000011101111100","001111010110110010100010010","001111010110001011000011010","001111010111100101100010100","001111010110100100011000010","001111010111110110001011111","001111010110010111100000001","001111010111110000010100100","001111011001001001110110111","001111011000011010100010001","001111011000010110111000010","001111011001000110101110001","001111011001000011011111100","001111011001011011101101111","001111010111001110111101100","001111010101011001111010100","001111010110111011100000111","001111010011110011000100101","001111010100010011000111101","001111010101010100101011000","001111010011000100010001111","001111010010111101011111110","001111010010001010000100010","001111001111110110010011001","001111010011010101011011110","001111010001101010101000001","001111010010111000110010111","001111010100100000011101001","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000"),
("000000000000000000000000000","000000000000000000000000000","001111010110111101000110101","001111010101111101100111011","001111010100010010101100011","001111010101010110000010000","001111010100011100010010111","001111010101000101101010100","001111010100010100100000110","001111010100000101101111000","001111010101001111101010001","001111010011010011000100110","001111010011101110001110010","001111010011010001000000101","001111010011101111011010110","001111010011100111011110010","001111010011011011010101010","001111010011110111000001011","001111010110001011000110011","001111010011111000111000111","001111010111101100100001001","001111010101000100101001100","001111010111011101111001111","001111010101010010001011101","001111011000010110101010101","001111011000000101101001110","001111011000000101010010101","001111010111011010100101000","001111010111000111111000101","001111011000011110000000111","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000"),
("000000000000000000000000000","000000000000000000000000000","001111010010010011100000010","001111001111110010001000111","001111010010000001000000011","001111010010010110000011111","001111010001110010101101000","001111010000101101001000110","001111010010000010111110010","001111010001110001100110110","001111001100111110110001000","001111001111110011101111101","001111001111111000110010101","001111010001010010101001000","001111001110010010001110100","001111010000000110000000110","001111010001100000111111100","001111010011011010011110110","001111010010111101100100000","001111010111011011001000101","001111010010011010101001100","001111010101010011110110100","001111010010111100111110010","001111011001000010111101000","001111010011111110001110110","001111010101010000110100101","001111010001110101100010011","001111010110011001000010101","001111010011101010010001100","001111010100010000000101101","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000"),
("000000000000000000000000000","000000000000000000000000000","001110111011111100100010110","001111001010111110000001011","001111001100101001111001001","001111010001000010001000000","001111010001111000001010010","001111010010110111010001010","001111010100101011010011011","001111010110000011101010010","001111011001000000000010111","001111011000100000001100111","001111011000011111111010101","001111011000000101110000100","001111010101111110101010100","001111010010110110000001101","001111001100100111000100110","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000"),
("000000000000000000000000000","000000000000000000000000000","001111011001000001010001000","001111010110110101110000111","001111010100111011110100010","001111010110101101000110001","001111010111000101111110111","001111010101010000001110111","001111011000011001111110100","001111011001111110101101001","001111011001000000110100001","001111010110000100010011010","001111010100111101010000101","001111010010111101001000110","001111010001000111101111101","001111000000100111000101111","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","001110111011101111111101011","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","001110111000011110001111101","001111001010000111000010010","001111001100111011011101010","001111001101101010011110101","001111010010011110010011010","001111001111000000001110111","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000"),
("000000000000000000000000000","000000000000000000000000000","001111010100101000110100000","001111010100100000110100010","001111010010101100101011111","001111010010111010000010100","001111010001100110001111000","001111010001101111110111101","001111010001000000011110001","001111010011000101100010101","001111010000011000101101010","001111001110010010101001110","001111001100100101110101001","001111001100101101001101000","001111001010001100011110011","001111001010101010000100001","001111001010010111011101000","001111001101010010100111111","001111010000111011111001100","001111010001011101001011010","001111010010001100001001100","001111010101000001100110011","001111010010010010100100100","001111010100111000010101000","001111010111001100000010111","001111010111110101101100011","001111011000000110111110001","001111010101101111100000100","001111011000001001100100111","001111010100101011111001001","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000"),
("000000000000000000000000000","000000000000000000000000000","001111000111000000111101000","001111000010110110101011100","001110111010100011000001010","001110110100001011000101111","001110101011000011110010011","001110100001100010010001010","000000000000000000000000000","000000000000000000000000000","001110001101111001001100010","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","001110111011010100010011011","001111000000111011001001010","001111000110101010011110011","001111001010010000010011110","001111001001000110000001100","001111001010001010011110100","001111001010101010000100001","001111001111000010011101100","001111001100100110010000011","001111001110110010011001111","001111001100100001101010110","001111001011000000101011010","001111001011001001110000001","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000"),
("000000000000000000000000000","000000000000000000000000000","001111010010110001100000010","001111001110010101000100111","001111001100101111010011001","001111001001101000100100000","001111001000111111100100011","001111000001011100101000101","001110111010010101010000100","001110111001111110101101101","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","001110110010010101011000111","001111001000001101110100111","001111010001000101000110111","001111010011000100111100111","001111011000101010011000001","001111011000110001111110001","001111011001101101101111010","001111011001011111011110000","001111011011100011000101010","001111011100101001000111111","001111011011101000100110000","001111011010110100111101100","001111011010100000110101110","001111011010010010110010001","001111011001010011100101110","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000"));
        wait for 300ns;
        wait;
        
    end process;
         

end Behavioral;
