----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 08.08.2023 11:18:39
-- Design Name: 
-- Module Name: fpupack - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;
package fpupack is
    constant FRAC_WIDTH : integer := 18;
    constant EXP_WIDTH : integer := 8;
    constant FP_WIDTH : integer:= FRAC_WIDTH+EXP_WIDTH+1;
    constant bias : std_logic_vector(EXP_WIDTH-1 downto 0) := "01111111";
    constant int_bias : integer := 127;
    constant int_alin : integer := 255;
    constant EXP_DF : std_logic_vector(EXP_WIDTH-1 downto 0) := "10000010";
    constant bias_MAX : std_logic_vector(EXP_WIDTH-1 downto 0) := "10000110";
    constant bias_MIN : std_logic_vector(EXP_WIDTH-1 downto 0) := "01110101";
    constant EXP_ONE: std_logic_vector(EXP_WIDTH-1 downto 0):= (others => '1');
    constant EXP_INF : std_logic_vector(EXP_WIDTH-1 downto 0) := "11111111";
    constant ZERO_V : std_logic_vector(FP_WIDTH-1 downto 0) := (others => '0');
   
    constant s_one : std_logic_vector(FP_WIDTH-1 downto 0) := "001111111000000000000000000";                                                               
    constant s_ten : std_logic_vector(FP_WIDTH-1 downto 0) := "010000010010000000000000000";                      
    constant s_twn : std_logic_vector(FP_WIDTH-1 downto 0) := "010000011010000000000000000";
    constant s_hundred : std_logic_vector(FP_WIDTH-1 downto 0) := "010000101100100000000000000";                                                                   
    constant s_pi2 : std_logic_vector(FP_WIDTH-1 downto 0) := "001111111100100100001111110";
    constant s_pi : std_logic_vector(FP_WIDTH-1 downto 0) := "010000000100100100001111110";
    constant s_3pi2 : std_logic_vector(FP_WIDTH-1 downto 0) := "010000001001011011001011111";
    constant s_2pi : std_logic_vector(FP_WIDTH-1 downto 0) := "010000001100100100001111110";
    
    constant Phyp : std_logic_vector(FP_WIDTH-1 downto 0) := "001111111001101001000001111";
    constant log2e : std_logic_vector(FP_WIDTH-1 downto 0) := "001111111011100010101010001";
    constant ilog2e : std_logic_vector(FP_WIDTH-1 downto 0) := "001111110011000101110010000";
    constant d_043 : std_logic_vector(FP_WIDTH-1 downto 0) :=  "001111010011000000100000110";
   
    constant MAX_ITER_CORDIC : std_logic_vector(4 downto 0):= "01111";
    constant MAX_POLY_MACKLR : std_logic_vector(3 downto 0):= "0011";
   
    constant OneM: std_logic_vector(FRAC_WIDTH downto 0) := "1000000000000000000";
    constant Zero: std_logic_vector(FP_WIDTH-1 downto 0) := (others => '0');
    constant Inf: std_logic_vector(FP_WIDTH-1 downto 0) := "011111111000000000000000000";
    constant NaN: std_logic_vector(FP_WIDTH-1 downto 0) := "011111111100000000000000000";
    constant TSed: POSITIVE := 15;
    constant Niter: POSITIVE := 3;
    
    -- PARAMETROS DA DIMEN?O DA CAMADA CONVOLUCIONAL
    constant sampleLength : integer := 66;
    constant inConvs : integer := 34;
    constant inConvs2 : integer := 32;
    constant outConvs : integer := 30;
    constant numberOfFilters : integer := 32;
    constant biasConvLength : integer := 32;
    
   -- ARRAYS PARA A PRIMEIRA CAMADA DE CONVOLU?O
    TYPE samples_adjust IS ARRAY ((sampleLength-1) downto 0) of std_logic_vector ((FP_WIDTH - 1) downto 0);
    TYPE filter IS ARRAY ((numberOfFilters-1) downto 0, 6 downto 0) of std_logic_vector ((FP_WIDTH-1) downto 0);
    TYPE biasConv IS ARRAY ((biasConvLength-1) downto 0) of std_logic_vector ((FP_WIDTH-1) downto 0);
    TYPE outConv IS ARRAY ((numberOfFilters-1) downto 0, 59 downto 0) of std_logic_vector ((FP_WIDTH-1) downto 0);
    -- ARRAYS PARA A SEGUNDA CAMADA DE CONVOLU?O
    TYPE in_Conv2 IS ARRAY ((numberOfFilters-1) downto 0, (inConvs-1) downto 0) of std_logic_vector ((FP_WIDTH-1) downto 0);
    TYPE filter2 IS ARRAY ((numberOfFilters-1) downto 0, (numberOfFilters-1) downto 0, 4 downto 0) of std_logic_vector ((FP_WIDTH-1) downto 0);
    TYPE aux_filter2 IS ARRAY ((numberOfFilters-1) downto 0, 4 downto 0) of std_logic_vector ((FP_WIDTH-1) downto 0);
    TYPE out_loop IS ARRAY ((numberOfFilters-1) downto 0) of std_logic_vector ((FP_WIDTH-1) downto 0);
    TYPE out_Conv2 IS ARRAY ((numberOfFilters-1) downto 0, (outConvs-1) downto 0) of std_logic_vector ((FP_WIDTH-1) downto 0);
    -- ARRAYS PARA A TERCEIRA CAMADA DE CONVOLU?O
    TYPE in_Conv3 IS ARRAY ((numberOfFilters-1) downto 0, (inConvs2-1) downto 0) of std_logic_vector ((FP_WIDTH-1) downto 0);
    TYPE filter3 IS ARRAY ((numberOfFilters-1) downto 0, (numberOfFilters-1) downto 0, 2 downto 0) of std_logic_vector ((FP_WIDTH-1) downto 0);
    TYPE aux_filter3 IS ARRAY ((numberOfFilters-1) downto 0, 2 downto 0) of std_logic_vector ((FP_WIDTH-1) downto 0);
     -- ARRAYS PARA A QUARTA CAMADA DE CONVOLU?O
    TYPE in_Conv4 IS ARRAY ((numberOfFilters-1) downto 0, (outConvs-1) downto 0) of std_logic_vector ((FP_WIDTH-1) downto 0);
    TYPE filter4 IS ARRAY ((numberOfFilters-1) downto 0, (numberOfFilters-1) downto 0) of std_logic_vector ((FP_WIDTH-1) downto 0);
    TYPE aux_filter4 IS ARRAY ((numberOfFilters-1) downto 0) of std_logic_vector ((FP_WIDTH-1) downto 0);
    -- CONSTANTES DOS FILTROS E BIAS ARMAZENADOS EM BROM DA FPGA
constant fourthConvBias : biasConv :=("001110101111011100001101101","001110111100000111011000000","001111001110110011010111010","001111010000101000001011000","101110111000100100000010110","001111001111110011100011111","001111001011010001111010110","001111001010101000100110011","001111001111001001001101101","001111001010110110110001110","001111001011101001110111011","001111000001111111101000010","001111010101000001100110111","001111001011001100111010001","101110111110000011011110011","001111010000001001100110111","001111001010101100110110000","101110111010010010000101101","001111001000101101010101000","001111001001100010100000110","001111011010011101111000000","001111000101010111110000110","001111000110001101010110110","001110111110110011001000001","001111001000011000010111110","000000000000000000000000000","001111010110101011010011110","101111000011011110101010001","001111010110011011101101101","001111000011101001011000111","001111010000101011110001011","001111000111010101100010101");

constant fourthConvfilter : filter4 :=((("101111100111101101100000110"),
("001111100000100110111011011"),
("101111011011110100101001001"),
("001111100001111101101110000"),
("001111100001101001010001011"),
("001111100000000100010010111"),
("001111100110111010001000100"),
("101111100110001111010111101"),
("101111101100100111011111001"),
("101111100000111010110001011"),
("101111101000101001010110101"),
("101111011011000010111000010"),
("001111010001110011101010110"),
("001111100100000001010110110"),
("001111100010000100110001001"),
("101111010110110000001000111"),
("101111011010011100111101001"),
("001111100100111101110001011"),
("101111100011010110110010101"),
("001111101011000100111000001"),
("101111011000111100011001111"),
("001111101000011110111010111"),
("101111101000100001010011110"),
("001111100000101100011010111"),
("001111011101100010101000110"),
("101111100110010100110110101"),
("001111101001010101110110100"),
("101111011100100001110100000"),
("001111100001001110000111111"),
("101111100110000100001100110"),
("001111100001110110000101101"),
("001111100001100000101101010")),
(("101111000010001011010111111"),
("101111011100010000101011010"),
("001111011000111100111100010"),
("001111101001010101100011001"),
("001111101000111100001100110"),
("001111100111001011010001110"),
("001111011011101011110111000"),
("001111100011110000001000001"),
("101111010111101101010100110"),
("001111011100010000110000101"),
("101111011011100000101110101"),
("101111101001001001101010010"),
("001111101001101001110100011"),
("001111100100001010010000001"),
("101111100110100100010011000"),
("001111100000011101111000101"),
("001111100110100111110101101"),
("101111100010100110101101111"),
("001111101010110110011001001"),
("001111010110101010101100001"),
("101111101000010000100001100"),
("101111101000010100100100010"),
("001111101010111110101110011"),
("001111101001000101001100010"),
("001111101001111000010011010"),
("101111101000110101111001111"),
("101111100010111101010000101"),
("001111101001100101000000000"),
("001111100011111011010111110"),
("001111010011001100110010100"),
("101111100001001100001011001"),
("101111011001000111011011111")),
(("101111011110010110100101100"),
("101111100101100101101010001"),
("001111001110110111010010011"),
("101111100101101000101101110"),
("001111010110001001011000000"),
("001111100110110100011101111"),
("001111101011000101111000011"),
("101111010011010101000010000"),
("101111011100011001001000111"),
("101111100110110101110010100"),
("101111001110101010110001001"),
("101111000001110001111011101"),
("101111100000001100000000110"),
("101111011101110110001111110"),
("001111100100100111001010000"),
("101111011111011111110011010"),
("001111100011001010000101100"),
("101111011111110100101000101"),
("001111010000001111011111000"),
("001111101011011101010100011"),
("101111011000001000110111010"),
("001111101001011101100111000"),
("101111100011011101000000001"),
("101111011000011001111101101"),
("001111100101111100000100101"),
("001111011111011111111001010"),
("101111100110011011110010011"),
("001111011001101001111110110"),
("001111011011011001110110000"),
("001111100110001110101011001"),
("001111001100101011111000110"),
("001111101010010100001011110")),
(("001111011110010100100101110"),
("001111101000111110111001111"),
("101111100100100010100101111"),
("101111010111100010101000011"),
("101111010110011110100011010"),
("101111010001110100000001111"),
("001111101011001111000000010"),
("001111010100101100000010001"),
("101111100111010110000010111"),
("101111010010111101001001000"),
("101111011011110011010011110"),
("101111101001010001011001011"),
("001111100001101101110001010"),
("001111011001001110110110011"),
("101111100111000010001101001"),
("101111011101001111110010011"),
("101111010111110001001111000"),
("001111011011010010001110101"),
("101111100110010001100001110"),
("001111100010111111101001111"),
("001111100000100010100110000"),
("001111101010011011100110100"),
("101111010000110000010101010"),
("101111101010101000110101101"),
("001111100111110101111010101"),
("101111100001111100010011001"),
("101111101001100101001010101"),
("101111100100110000100101111"),
("001111011010001011010010110"),
("001111100001110100010011010"),
("001111101000010101100111010"),
("001111011100001010000100111")),
(("101111100111001110110100110"),
("001111101001010001010001000"),
("001111011111011001011110001"),
("001111011110110011101010101"),
("001111011100100000011000010"),
("001111011111101100000110100"),
("001111100001010000111100100"),
("101111011111011101111100100"),
("001111011001000001010001101"),
("001111100111111011100000110"),
("001111100000100111111010111"),
("101111101010011001011011111"),
("001111010110011010101101110"),
("001111011011010101000011010"),
("101111001001101010010000110"),
("101111100111011111111100111"),
("101111000100110001011011100"),
("001111011111000100100100111"),
("001111010111100100001101111"),
("001111100010101101000110111"),
("101111101100100100011100000"),
("001111100000111101000000101"),
("001111101001000010110101001"),
("101111100111000100111100010"),
("001111101011001110101111101"),
("001111100111110110000111000"),
("001111010011110010011101001"),
("101111100010100111001101111"),
("101111100000111100001011010"),
("001111100111011011110000001"),
("001110111001000011001100000"),
("101111101000101110010101110")),
(("001111100110100000111110011"),
("001111101001010101010111011"),
("101111100100100110001011011"),
("101111011000011001100000110"),
("101111100101010111001010001"),
("101111101001110010010111001"),
("001111101000001001011011011"),
("001111011101010100010000001"),
("001111001000010101110101010"),
("001111100010100000101000110"),
("101111101000100010110001010"),
("001111011100000110101011010"),
("001111100110111010100110100"),
("001111100110010110110011110"),
("001111100100011010001100110"),
("101111100011000010110100010"),
("101111010101010001001010001"),
("101111000101111101000100111"),
("001111101000101000010110101"),
("101111100100110100110010100"),
("101111011001001100010111001"),
("001111001100011111110111010"),
("001111011011011011100111110"),
("001111101000011101010011000"),
("101111011011100010011000111"),
("101111100100111101000100000"),
("101111100011001000010010001"),
("001111100111010110010110111"),
("001111011000101000111111111"),
("101111100010111110111000010"),
("101111100111011110001110010"),
("001111011110000111100000111")),
(("001111100001010000001000001"),
("101111011010011110110111000"),
("001111100010010000111101010"),
("101111010001111101010111001"),
("101111011111111011000000000"),
("001111101010110011100100000"),
("001111100000110100000001100"),
("101111010101001101101111101"),
("101111101011110001101110010"),
("101111000000001000000011010"),
("001111100001111101001001101"),
("001110100000011111000010010"),
("101111010010111001110001010"),
("001111100110001010010000111"),
("101111100111101000111010001"),
("001111101000010000010101101"),
("001111000010010110010100011"),
("101111011000010110100000010"),
("001111100011000100100000000"),
("001111100111111111101101011"),
("101111011000110111100111101"),
("101111100001011011001100000"),
("101111011001110101011101010"),
("001111100001110001100010111"),
("101111101001000100101000111"),
("101111011111001001111001010"),
("001111100010111001111111011"),
("001111100011001111010011010"),
("101111100100111000111010101"),
("101111100001001110010000001"),
("101111100111101100010010001"),
("001111101010100010110001000")),
(("101111100000111101101110001"),
("001111100101010101111111100"),
("101111101010100100011010001"),
("001111100001000101101101110"),
("001111010001010110110101001"),
("001111011011000100001011000"),
("001111100011110001110110001"),
("001111011011001110000001010"),
("101111100000000110110001010"),
("001111100101110111001000011"),
("101111100011100001100110010"),
("101111100001001000100111111"),
("001111001101010101001001010"),
("001111100110100001011001011"),
("001111011110011111010011101"),
("001110010001000110101000000"),
("001111100010010111001110100"),
("001111011101100011100100010"),
("001111011100000000100111010"),
("001111100101010001110100101"),
("101111101010111001100101111"),
("001111000111000110110110101"),
("101111011110111101010111010"),
("101111100101101111000000110"),
("001111100001011111101010000"),
("001111011010001000101001111"),
("101111011001010000111111110"),
("001111011010000000000110000"),
("001111100111010000110000110"),
("101111001000101110100001011"),
("101111100111100001111000101"),
("001111101000100110011000001")),
(("101111011001011011101101101"),
("001111011000010000101000010"),
("001111100011010010110101000"),
("001111011000110111110011110"),
("101111010100011110111011110"),
("001111011111010001110100001"),
("001111100101011100110110011"),
("101111101001101010100001010"),
("001111100100001011101111111"),
("101111100011011011010111100"),
("001111100111111100001010001"),
("001111100011111101000100011"),
("101111001110000001001001000"),
("101111010100110111100100000"),
("101111011011111101101011010"),
("101111101000011101010100110"),
("101111011000101010111111111"),
("001111011111000010101100000"),
("101111101001000100101001110"),
("001111101000010111100111111"),
("101111101000100100111010111"),
("001111100000011000100100111"),
("101111100110011101010001110"),
("101111100011011010101001101"),
("101111100011101111001001011"),
("101111101000100101101000111"),
("001110111000011101001010110"),
("001111101001000001100011011"),
("101111100011000000001111000"),
("001111101001011010100101110"),
("101111011110100001111111111"),
("001111101001010100000000111")),
(("001111001011000101100100110"),
("101111100001111100100110001"),
("001111100011111110010000101"),
("101111010111011110001110001"),
("001111100100100011101111010"),
("001111101011001000010011100"),
("101111000000111111100001011"),
("101111100100000001011100100"),
("101111011100100000001101110"),
("001111100100001100000010101"),
("001111100001111101101001010"),
("101111101010100000011111100"),
("101111101001000010000010100"),
("101111011011111110011100111"),
("001111100110011011011000111"),
("001111101000001000111101001"),
("001111001011011101110100010"),
("001111001110001000011110010"),
("001111011011000011111101100"),
("001111011110101100101011100"),
("101111100100100000001010001"),
("101111000111110101100111010"),
("001111100000111110110100110"),
("101111101000000001111101010"),
("101111000100101010111101101"),
("001111100001011100011101110"),
("001111101000110011001000011"),
("101111100000010110000101011"),
("001111101001001010110001100"),
("001111101001100001111110001"),
("001111100001010010000101001"),
("101111011011001101110111100")),
(("101111101000000010000010001"),
("001111101001000111110101001"),
("001111011000011000001111000"),
("101111100011001000100110110"),
("001111001000111000001110011"),
("001111011100111001100010000"),
("101111011101111110000100001"),
("001111100000001111101011000"),
("001111101001011000101111100"),
("001111100011111011000110111"),
("001111001000100011111101001"),
("101111011001101101111001001"),
("001111011011101010001101111"),
("001111100011001101000011011"),
("001111100001111010101111000"),
("001111100010110000011000111"),
("001111101000011001001111100"),
("001111000000011111010100001"),
("101111101000001000110011110"),
("101111100010101111010110100"),
("001111011010001110100100010"),
("101111000010010001010101010"),
("001111101000010010101110110"),
("001111100100011110111010111"),
("001111011110010011101000001"),
("001111101000001100100110110"),
("001111100011111011011100110"),
("001111010011110010001011000"),
("101111100001001111010100011"),
("001111101000110101000010011"),
("001111100101100000001000010"),
("101111100111010001111001111")),
(("001111100101010001110011101"),
("101111100011111010110101010"),
("101111010110110001110110100"),
("001111100101010101101001011"),
("001111001101111110101101001"),
("001111100001000111100001011"),
("001111101001110000110101000"),
("101111101000101110101010010"),
("101111000010010110101010001"),
("101111100000011010001000101"),
("001111100010000111010000110"),
("101111010011111100110111011"),
("101111100110101110000001000"),
("101111100011000000110001101"),
("001111010010101011000100011"),
("001111011101001110000110100"),
("001111100001010000110101000"),
("001111100111010001100110101"),
("001111100111101110101110100"),
("001111100000010100111100000"),
("101111100010000011101110100"),
("101111100011001111111100011"),
("001110111011010110101110011"),
("001111011100010101100101100"),
("001111101001001110000011101"),
("001111101001111110001110110"),
("001111101010011000100110111"),
("101110111001111010111011111"),
("001111101000011111110100010"),
("001111101001011100100111010"),
("001111011100011011010110101"),
("001111100100000100010110000")),
(("001111000001101110100001110"),
("001111101000111001011001001"),
("001111011000011110000111111"),
("101111100001100111111000110"),
("101111100101011111110110001"),
("001111011101001011010000110"),
("001111101010011110001101001"),
("101111010000010001000100011"),
("101111100010011100101110111"),
("101111100101100100011011110"),
("101111011010100110110001101"),
("001111100001101100001101010"),
("001111101001001110111110111"),
("001111100110101111111100000"),
("101111101000101001000100001"),
("101111011110010101011111000"),
("101111011100010100001111010"),
("101111010001001011011100101"),
("101111011110010011110100010"),
("101111010111000001011110100"),
("001111011110111001000000111"),
("001111100011000100111011011"),
("001111100011100101001101001"),
("101111100100010000001010010"),
("101111101010010010001011011"),
("101111100100011111110001001"),
("101111011011110101001011101"),
("001111001010101010011010110"),
("101111100011001000000010110"),
("001111100001000100000011111"),
("101111101001110110100111011"),
("001111101010010111100011111")),
(("001111100000110110111101010"),
("101111100011001111100101011"),
("101111101011010001010000000"),
("001111101001010000010111110"),
("101111011110011001010110111"),
("101111000101100011110110000"),
("001111100010000000001001011"),
("001111100010001011101011000"),
("001111100101101111100000100"),
("001111001011000100001101010"),
("101111100101010000101101010"),
("101111010111001010110111110"),
("001111011010101000100001001"),
("001111100110011110001010101"),
("001110110110010000001001110"),
("101111100111101111101010100"),
("101111100110011010010001011"),
("101111001110110101100001011"),
("001111100010000111011110100"),
("001111010111001011011011011"),
("101111011100000100010001000"),
("001111011011001011110001010"),
("101111100100111010100100111"),
("001111010001111100110110100"),
("001111010010011100100100011"),
("101111100001011000000110110"),
("101110010001111110101111111"),
("101111011111111001111101010"),
("101111100100110110101100111"),
("101111101001001011000001001"),
("101111100011011100010111101"),
("101111100001011000011011111")),
(("101111011010101111010001111"),
("101111101001101010011001011"),
("101111100101001101110111001"),
("001111011101110100100110010"),
("101111101000011100100111101"),
("001111011010110101001001000"),
("001111011000000100000111000"),
("101111100101100110000110000"),
("001111011110011111100010101"),
("001111011110110110001100110"),
("001111100101001101001010010"),
("001111100010001111000100001"),
("101111000101001010010011000"),
("101111011011100010100001000"),
("001111101000010001000100001"),
("001111011111101001111110101"),
("001111100011110001000111001"),
("001111101000111101000110101"),
("101110100101111101110101100"),
("001111010011010111000110011"),
("101111100001001110100001011"),
("001111100010100001001100000"),
("001111101010000011111011100"),
("001111011111011110000101100"),
("001111010110011010011001100"),
("001111100000111110001111101"),
("001111100101011000110111010"),
("001111101010010101000011010"),
("101111100011110011000100111"),
("101111100000100110100101001"),
("101111100101010011111010110"),
("001111100000010110101110111")),
(("101111101000110010000101000"),
("001111010101101011000010101"),
("101111100011001110000010000"),
("101111010011110001000010111"),
("001111100101010011100100001"),
("101111101010011011110001100"),
("001111101011001101010110111"),
("001111100011001110001101110"),
("101111001001011011110011010"),
("001111101000001011110001000"),
("001111101000010100000000000"),
("001111001010110111100001100"),
("001111100000000101111110101"),
("001111100110101110101000011"),
("101111101001011101111000001"),
("101111011000100001101011000"),
("101111011110111101010011100"),
("001111100000100101101110101"),
("001111100110000010111110110"),
("101111000101011010000010110"),
("001111010010111100110011000"),
("101111101001001011001011111"),
("101111101000000111111010000"),
("001111101001011001100100010"),
("101111101001011101011101011"),
("001111100011010110000011000"),
("001111101000110011100000001"),
("001111011011101101010100100"),
("101111011100010100010011111"),
("101111100100011101100001000"),
("001111001111100010011110000"),
("001111011000100001000000101")),
(("001111100111010011010010100"),
("101111101000111011110001111"),
("001111011100001110011111100"),
("101111101000001001100100100"),
("101111100000011100011011100"),
("101111011111101110001100111"),
("101111011010011010010010100"),
("001111100010111001111011010"),
("101111011001011111101110111"),
("101111101000010100101000111"),
("101111100111100011100111000"),
("101111101001000111110000101"),
("001111011101001110011100000"),
("101111100001110000000110011"),
("001111101001110010001101011"),
("101111001011100000001011000"),
("001111100010101110111011000"),
("101111010001111011011101001"),
("101111100010100100000111001"),
("101111101001001000111110101"),
("001111011000011010100111010"),
("101111011011110110110100000"),
("001111011010011001100001101"),
("001111011010101110011110111"),
("101111101010110001001100001"),
("101111011000000100101000111"),
("001111100001011100100001101"),
("101111001011010101001111100"),
("001110101011000111000001111"),
("001111100001001101101000100"),
("101111101001000001001000101"),
("001111101001001010111111000")),
(("101111011010000000000110110"),
("001111011111100110110011100"),
("001111100111010011010010101"),
("101111100110010011100101101"),
("101111100100110010100110000"),
("001111010000100001011111000"),
("101111100010001000101110001"),
("001111011001101001101001100"),
("001111100001010001100010010"),
("101111100000101101010100010"),
("101111101010110010011001001"),
("101111100001010111101010001"),
("001111100100000001111101111"),
("001111011010010100110000110"),
("001111011100110100101101000"),
("101111100101111000101011000"),
("001111100100001011111001010"),
("101111100001000010111101111"),
("001111101001011011111011110"),
("101111100100010001011010110"),
("001111101000000101110111100"),
("001111100000000000001000011"),
("101110111010100110110010000"),
("001111100101000000100001001"),
("001111100111111001001000110"),
("101111100000110011110010001"),
("001111001001010010011010000"),
("101111101000000010111101110"),
("001111100111001001011101100"),
("101111011111010110101100111"),
("001111000001111000011100000"),
("001111100111111010010100011")),
(("001111101001000110110011101"),
("001111100100101010101100100"),
("101111100010111111011111001"),
("101111100000100111010101011"),
("001111100101110000111011010"),
("101111010110001100101011001"),
("001111001111011101001111000"),
("101111010000111000110001010"),
("001111011011111001100110010"),
("001111011110110110010011000"),
("001111100100110010100100111"),
("001111010001001000001111101"),
("001111001000101000111110000"),
("001111101000110010110110000"),
("001111101000110010100110110"),
("001111101001011000101010110"),
("101111100000111001000110101"),
("101111100011101001001111110"),
("001111010001111111111100000"),
("101111100111011110011010010"),
("101111101000011111010001011"),
("001111100111001010100110000"),
("001111100010110011110000111"),
("001111100011010010110100110"),
("101111011110001110011110111"),
("101111101000010110111011100"),
("101111011010000101000101110"),
("101111101001011001101011110"),
("101111100100011000111011111"),
("101111011001011111100000100"),
("101111001111110111010011100"),
("101111100011100010110101011")),
(("001111100111101000110010000"),
("101111101001101110000001100"),
("001111010010111100111101110"),
("101111100111010100101010000"),
("101111001001101101111111110"),
("101111100011111001110100001"),
("001111101001111111100111010"),
("001111100101000001000001110"),
("101111101000111100111000111"),
("101111101000101010101011100"),
("001111101001101010001000010"),
("101111100110100001101111010"),
("101111100111011111110101011"),
("101111010110101001101010010"),
("101111100000000001111010110"),
("001111010110010101101111100"),
("001111001000110111111010100"),
("001111100000001010100011011"),
("101111011110100100010010111"),
("101111011010111001000100001"),
("101111011100010100110000101"),
("101110111101111010001111000"),
("001111011101010100010011110"),
("101111100101000110011111001"),
("001111000001001100101101111"),
("001111011011011000000110000"),
("001111101000111011000110000"),
("101111100101011100101010011"),
("001111100101000001111100010"),
("001111100101011001001010101"),
("101111100000111110001100111"),
("001111100011111000100100101")),
(("101111000110001010111000111"),
("001111011110011011011010000"),
("101111010011111110000011111"),
("001111100101111010001110111"),
("001111100011101010100000011"),
("101111101000010010001011111"),
("001111100111001010011100111"),
("101111100000000111101110001"),
("101111101010010101001011000"),
("101111010100010111000010011"),
("001111010001110010000010111"),
("101111011000010100101101111"),
("001111100100010100110000110"),
("001110110010011110010010100"),
("001111010110000010110111000"),
("001111100101111111001001100"),
("101111100011011010100011011"),
("001111101010101100011010000"),
("101111100101100100110111011"),
("001111000101101010100100010"),
("001111101001101101111011001"),
("101111011000010010111101011"),
("101110110110011111100111111"),
("101111100100110011110110010"),
("001111100101010100111011101"),
("001111011101100011001000000"),
("101111001010110001101001111"),
("101111011000010110101111111"),
("101111101000110110000010000"),
("101111100111100001101110001"),
("001111001000110001010101100"),
("101111100001100010010010110")),
(("001111101011001000101100101"),
("001111100101101111010011100"),
("001111011010000000110001111"),
("101110110111011010110100010"),
("101111100001100111100000000"),
("101111101000101111111010111"),
("101111011110111100000100100"),
("101111100011111010010110000"),
("001111101000001011111110111"),
("001111100100011101011000011"),
("101111100001011110101000100"),
("101111100111101110010110100"),
("001111100010011011110010010"),
("001111100000001001000011000"),
("101111010110010111110100101"),
("001111100110101011111100110"),
("101111011100110000101110111"),
("101110100001100101011111100"),
("001111010010100011001111110"),
("001111010111000001100110010"),
("101111011011100101000101010"),
("001111100010111101000111011"),
("101111100011110010000101011"),
("101111100101110001011111011"),
("101111101001100010000101111"),
("101111011001101100101001100"),
("001111100111100010100101001"),
("001111001011011011111110111"),
("101111100010100011101011101"),
("101111100010000001111111001"),
("101111101001100011000001001"),
("101111100011100000111011101")),
(("101111101000010111110011001"),
("101111010010010111110000000"),
("101111100101000111111010110"),
("101111010101110011000101010"),
("101111011000010011001000010"),
("001111101001000000001111110"),
("101111100100000001010100010"),
("001111100100101010010100000"),
("001111000001100110010000100"),
("001111100010011100101110010"),
("101111101000011011110101011"),
("001111100000111010111111011"),
("101111100000011010110101010"),
("101111100000110110100010010"),
("001111100011110110001100110"),
("001111100110101000011010010"),
("001111100101111000000100000"),
("001111101010111100011011000"),
("001111011001000001110000001"),
("001111101010001000010010101"),
("001111100110010011011100000"),
("101111100011011101000101010"),
("001111001110010111111011110"),
("101111100001000110011000101"),
("101111100001100111100101100"),
("101111100000100001100110001"),
("001111100011000101011010010"),
("001111101011101111100111110"),
("101111100011011001010101001"),
("001111100111100011011110101"),
("001111100100010000101001010"),
("101111101001100011001011000")),
(("001111101000101011101101000"),
("101111001000010101000101100"),
("101111100100100001011010001"),
("101111101001010111001101011"),
("001111101001110010100010001"),
("101111100100100101001111000"),
("001111011011110111001101000"),
("101111001011000110110111101"),
("001111100001101111000010010"),
("001111011100011111100111111"),
("101111100001101001010001001"),
("001111101010010010110011000"),
("101111010101001001111010110"),
("001111011001110100001001111"),
("101111010110010000010010010"),
("001111000110001110111100110"),
("001111100101000011000011111"),
("001111101000100110011000011"),
("001111101000100110100001011"),
("001111010011110110110100101"),
("101111011010001100101110010"),
("001111100111100011111101010"),
("101111100101111010011001010"),
("001111011001001000001000101"),
("101111101000101110101000000"),
("101111101010100001100011000"),
("101111100101001001011011111"),
("101111101010001010001011111"),
("001111100000010110100000000"),
("101111011010010010011100110"),
("001111000111111001001000011"),
("001111101010100100001011000")),
(("001111101000000000110001010"),
("001111100111111010011011111"),
("101111100111100111001111000"),
("101111010000110011100101010"),
("001111011011000100110100100"),
("101111001000001010001000100"),
("001111100010011000111100010"),
("101111010110100001110100010"),
("101111011101110111110110010"),
("101111101001010110100010011"),
("001111101001101000001111110"),
("001111100000011010010110010"),
("001111011011110001101111100"),
("001111100011011111101100100"),
("001111100011101011111010101"),
("001111010011000010001100001"),
("001111101000000111100101001"),
("001111011111000100110011110"),
("101111101011110110100001110"),
("001111101011000011011101000"),
("001111010010111011101000000"),
("101111100010100000110110100"),
("001111100101010111100000100"),
("101111100101011001111101011"),
("001111010000001100010010011"),
("101110100100001110100010100"),
("101111101000010000101001100"),
("101111011101110010010011000"),
("101111100101100110100000010"),
("001111100010100110001101110"),
("001111101000110101101010111"),
("001111100001000111010001010")),
(("001111010001101000011000011"),
("101111100011001010011001011"),
("001111100011001010111110111"),
("101111011000111001011101110"),
("101111100111110010110110101"),
("101111100000111000011000100"),
("101111100110011100001111000"),
("101111101000001101001111011"),
("101111101000110010010110011"),
("101111100100110011101010010"),
("001111100010001100101100100"),
("001111011001110011101010000"),
("001111101000101011011110101"),
("101111101000001100100111100"),
("101111100111011100010010101"),
("001111100111001001110000010"),
("101111101001101000001001101"),
("101111011110110011100010101"),
("001111100110001001111010001"),
("001111100111001101111010001"),
("101111100010011101001101101"),
("101111010011111010100000011"),
("101111100101001101100001010"),
("101111100101101001011111100"),
("101111010101010111010110001"),
("001111001111010111011001000"),
("101111100000111000111100011"),
("101111101000100110101001011"),
("101111011001101101110111110"),
("001110101101011010111001000"),
("101111100101110100000011110"),
("001111010010010001100001100")),
(("001111101001000100010010000"),
("001111000001000111111110110"),
("001111101000111100010100101"),
("101111100101011111100111111"),
("001111101001101001110001001"),
("001111100100110101111111010"),
("101111010000000011000100011"),
("001111010111000110111010100"),
("101111101010000010101011001"),
("101111011110100011001101110"),
("001111100110000101011011010"),
("101111100000100111111001101"),
("101111100001110110011101010"),
("001111100101000001011011110"),
("101111010111111111011100001"),
("101111011100100100001110100"),
("101111100000000101011001111"),
("101111011110110110000011001"),
("001111010101110010100001100"),
("001111101000111100110000000"),
("001111101001100000000110111"),
("001111100000001011011001000"),
("101111100100111111001001001"),
("101111100001101111111000010"),
("101111010111001000001000111"),
("101111100010100000011010000"),
("101111100110110001011100111"),
("101111011111000100101001001"),
("101111101000001010111001100"),
("101110110111100010000010110"),
("101111101000001110100010001"),
("001111101001100111101010001")),
(("101111100100101010000101101"),
("001111100000111001011100111"),
("101111100000111011111011001"),
("101111101001001010001111011"),
("001111010011100111010111110"),
("101111100001110000110011011"),
("001111100101001111010011001"),
("001111011101001111001011100"),
("001111011110111100010110010"),
("001111011011001001101010000"),
("101111011100101011000110000"),
("101111100011001111100011101"),
("001111011110000110100101010"),
("101111100011010001011001000"),
("101111011001111010000111110"),
("101111101000000010110000000"),
("101111101000011101001100000"),
("001111100010101001100100110"),
("101111101000001000101011111"),
("101111101001111010100010111"),
("001111101010010000011111110"),
("001111100010011100000110101"),
("101111010110001010101001111"),
("001111101001010101000110000"),
("101111001000000101001000011"),
("101111011110100111010010010"),
("001111100111100011100000110"),
("001111101000110010110100111"),
("101111101010111100001010110"),
("001111101001111111011010100"),
("001111011011100011000110010"),
("101111001101011110110001111")),
(("001111100101011110110111010"),
("001111100100101001110101000"),
("101111011101110001110100001"),
("001111100100011100100001011"),
("001111011000001001110111101"),
("101111100100101111101010011"),
("101111011101000110100001011"),
("001111101000101011010011000"),
("101111100011110000011110001"),
("001111101000101010100010101"),
("101111011010101100000100011"),
("101111100111010101011110100"),
("101111100111010110011001110"),
("001111101001000111000011100"),
("101111101000000111010101000"),
("101111010010101010100110111"),
("101110110101000010011100100"),
("001111001100111111000001000"),
("101111100100111100011111000"),
("101111010101001010000010010"),
("101111100101000111011010111"),
("101111100000100011100011110"),
("001111011010111000010011011"),
("101111011011100100010010011"),
("101111101011111000101101111"),
("001111100110100100001111110"),
("101111101001100010100110000"),
("101111101000001110000011101"),
("001111101011001010001011110"),
("101111100010110110100000101"),
("101111100011010111111011010"),
("001111101001011101011011000")),
(("101111100010111110011111110"),
("001111011101010000000101010"),
("001111101001111101100101010"),
("101111101000010100111001111"),
("101111000011001010010100010"),
("001111101000000001011010001"),
("101111100111101110100111010"),
("001111010111010000100000001"),
("001111100011001101111010101"),
("101111001111100010100011000"),
("101111101000000000111101001"),
("001111100100100001110101000"),
("101111100000111110101111100"),
("001111001011010000100100011"),
("001111000110010011110111000"),
("101111100010000000010101011"),
("101111100101000001011100100"),
("001111100101010010111010001"),
("001111101000010010100111110"),
("001111100011001101001100100"),
("001111010110001001111000010"),
("001111101000001110001101111"),
("101111100100000111011011000"),
("001111100101011111111010011"),
("101111101000110000010010110"),
("101111100100100110000110101"),
("001111101001110001100101001"),
("001111010001101101011110000"),
("101111101001101100101000101"),
("001111101010000100000001001"),
("101111100011101011110101100"),
("101111101001010110010111001")),
(("001111101001110010000001011"),
("101111100000010100010010100"),
("001111011111100010011001000"),
("101111011100011110110100001"),
("101111010001010111101001001"),
("101111011010100010011111110"),
("001111100010011011010001010"),
("001111100100001011111100010"),
("101111100100001000110011000"),
("001111010110000000010110111"),
("001111011100100111110011110"),
("101111010000010101101111101"),
("001111001110101100011110111"),
("101111100101101001101100001"),
("101111100110010001101110110"),
("101111101000001110010110011"),
("101111100011110010000010110"),
("101111100000011011011011000"),
("101111100010100000000101001"),
("001111100110110101100111110"),
("101111100111101010111001101"),
("001111011101011100011011010"),
("101111100000000010001000000"),
("101111011110111111011000011"),
("001111100110100000000000110"),
("101111100101110001111001000"),
("001111011110110100000010001"),
("001111101001100001110110101"),
("101111100010001110110110100"),
("001111101000100110110100111"),
("001111100110111101011010011"),
("001111100011000100000001010")),
(("001111100111010100001001000"),
("001111101100011001111101000"),
("101111100010110111010010000"),
("001111100000110010010100111"),
("001111101001001011010011101"),
("001111011111001000101011000"),
("001111011000110011010100010"),
("001111100110111001000001001"),
("001111101000001101010000101"),
("101111101001001100101100101"),
("001111101011111100101011001"),
("001111011001010011000111110"),
("001111101000010101000000010"),
("001111011100001000000010101"),
("101111101000110101010110110"),
("001111100101010101110110011"),
("101111011111000000100101001"),
("101111010010101000011100000"),
("101111011111000111101001101"),
("001111101010001111001001000"),
("001111101000010111010111111"),
("101111100001000000010101001"),
("101111101001000010101010100"),
("101111011110010000001010110"),
("101111011000011000001100000"),
("101111100001000101111010001"),
("101111101001111001111101111"),
("101111001011001110011100100"),
("101111101010101000001101101"),
("001111010010101100111010001"),
("101111100011110111010111111"),
("101111100111101011001001011")));
end fpupack;

package body fpupack is
end fpupack;