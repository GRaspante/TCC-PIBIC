----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 07.08.2023 21:29:38
-- Design Name: 
-- Module Name: cnn_conv3c_tb - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_unsigned.all;
use IEEE.NUMERIC_STD.ALL;
use work.fpupack.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity cnn_conv3c_tb is
--  Port ( );
end cnn_conv3c_tb;

architecture Behavioral of cnn_conv3c_tb is

component cnn_conv3c is
    Port (   reset_conv3 : in STD_LOGIC;
            clk : in STD_LOGIC;
            start_conv3 : in STD_LOGIC;
            samples_conv3 : in in_Conv3;
--            filter_conv3 : in filter3;
 --           bias_conv3 : in biasConv;
            ready_conv3: out STD_LOGIC;            
            out_conv3: out std_logic_vector (FP_WIDTH-1 downto 0));
end component;

signal sreset_conv3, sclk, s_start_conv3, sready_conv3 : std_logic;
signal s_samples_conv3 : in_Conv3;
signal sfilter_conv3 : filter3;
signal sbias_conv3 : biasConv;
signal s_out_conv3tb: std_logic_vector (FP_WIDTH-1 downto 0);

begin
uut: cnn_conv3c port map (     reset_conv3       => sreset_conv3,
                                clk               => sclk,
                                start_conv3       => s_start_conv3,
                                ready_conv3       => sready_conv3,
                                samples_conv3     => s_samples_conv3,                                    
                           --     filter_conv3      => sfilter_conv3,                                
                          --      bias_conv3        => sbias_conv3,                                
                                out_conv3      => s_out_conv3tb);
                                
clk: process
        begin
            sclk <= '0';
            wait for 5ns;
            sclk <= '1';
            wait for 5ns;            
        end process;
        
stimulus: process
    begin
        sreset_conv3 <= '0';
        s_start_conv3 <= '0';            
        wait for 10ns;            
        sreset_conv3 <= '1';
        s_samples_conv3 <= ((others =>(others => (others => '0'))));
        sbias_conv3<= (others => (others => '0'));
        sfilter_conv3 <= ((others =>(others =>(others => (others => '0')))));
        wait for 20ns;
        
        sreset_conv3 <= '0';
        wait for 10ns;
        
        s_start_conv3 <= '1'; 
        sbias_conv3 <= thirdConvBias;
        sfilter_conv3 <= thirdConvfilter;
        s_samples_conv3 <= (("000000000000000000000000000","001111001111101000000101000","001111011000000001001000010","001111011011011011111001111","001111011100111011101101000","001111011110011010000000000","001111100000001111000000001","001111100000111110101111110","001111100001100100100110100","001111100010000101100010111","001111100010010100101110011","001111100001011001011000100","001111100000001000010111100","001111011100100011100001110","001111011000001011100101110","001111001111010110010110100","001110110010101001000011001","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","001110111101010001110111101","000000000000000000000000000","000000000000000000000000000"),
                        ("000000000000000000000000000","001111001011000010000011010","001111001100011111011000000","001111010111001011010011110","001111010111000101000111011","001111010100110100001000100","001111010111011100000010011","001111011000111000111101111","001111011010000011111011101","001111011010011111001110100","001111011010100001110011101","001111011001110001011110011","001111011000010110011100100","001111010100101011011011110","001111001101110000000001000","001111000000101101100101001","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","001111000001111010001000000","001110111111110001101001011","000000000000000000000000000","000000000000000000000000000"),
                        ("000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","001110110111101001011000111","001111001100110000001101111","001111010010000010001111001","001111010001011111111010010","001111001110001001011000010","001110111111101100100010010","001110111111101011101111111","001110101010010110101100110","001111000100011011100010101","001111001010000010101001010","001111001010111000001110001","001111010001011010001010010","001111010001100010000011101","001111010011111101010001111","001111010001011100100101100","001111010011001010011000000","001111010001010100100101110","001111010011110110010110011","000000000000000000000000000","000000000000000000000000000"),
                        ("000000000000000000000000000","001111100001000110000101010","001111100100011100100000100","001111100101100001011010100","001111100100110100001000000","001111100101011101101010101","001111100101111110110000100","001111100110010111011101110","001111100110000000100011101","001111100110000000001000101","001111100100100010000011011","001111100011001000011100000","001111100000111001000010100","001111011110100101110110001","001111011011010011010101100","001111011000111100000100000","001111010010111001011111111","001111010011010010100110011","001111001110000010011011101","001111000111111000000000010","001110101001111000110100001","000000000000000000000000000","001110110010110011010001100","001111001011111110111011110","001111010111010101100110010","001111011011110000100000000","001111011110001100110011111","001111100000010000010110001","001111100001100111001101001","001111100000011010111001011","000000000000000000000000000","000000000000000000000000000"),
                        ("000000000000000000000000000","001111100010100000001111110","001111100100100010010010111","001111100101111111010010000","001111100101100111011011011","001111100101010111010010010","001111100101101000010100100","001111100101100101011001010","001111100101001110100100111","001111100100001111100010100","001111100011011100010001000","001111100010110111110101010","001111100010010000101010001","001111100001010100111110101","001111100000110010101001011","001111100000110001000001010","001111100000101110111010100","001111100000001111001001001","001111011100110100100111100","001111011001100000010111001","001111010010111011011101110","001111000101001110110010100","001111000010010001011101010","001111010000000101111000011","001111010100010011101000001","001111011010110010000111000","001111011110111010110000101","001111100001111000110010000","001111100011100001111110001","001111100011001111000000110","000000000000000000000000000","000000000000000000000000000"),
                        ("000000000000000000000000000","001111001011000110111001101","001111010100001011000101111","001111011001111001101110111","001111011001001000100111010","001111011001010010111110100","001111011010000000110000001","001111011010111000001100000","001111011010010010000110101","001111011001111110101111010","001111011001001010011010000","001111010101000011011111000","001111010001001100000001011","001111001001000110110110000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","001111001011011100110000100","001111010000110001110101110","001111001111011100010000000","000000000000000000000000000","000000000000000000000000000"),
                        ("000000000000000000000000000","001111100010001111010010100","001111100100000110000101100","001111100101010100010010011","001111100100101010110010010","001111100100011001011100011","001111100011111110011111110","001111100011100011111111011","001111100011010010010011110","001111100011010100110111100","001111100011011110110100111","001111100011001001010000101","001111100011010100000111011","001111100011100010010011011","001111100011101111011110100","001111100011111001101010111","001111100011001010000100100","001111100001111110100110100","001111100000001011001111110","001111011011001111011110101","001111011001010001100010110","001111010100000101110001000","001111001111010100100001000","001111001111111110011111100","001111011000001111000000011","001111011100101101110100010","001111011111000111010011011","001111100010011000111001100","001111100010110101000001011","001111100010000000001010101","000000000000000000000000000","000000000000000000000000000"),
                        ("000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000"),
                        ("000000000000000000000000000","001111010111000101000011001","001111011011001000011010101","001111011010110010110111010","001111011011010001110011000","001111011011010100111011010","001111011011101000011011100","001111011011110111010010001","001111011100110000011110101","001111011110101001101100101","001111011110001101101001011","001111011110101111101110100","001111100000000100110000110","001111100000001100101000101","001111100000000011100110001","001111011110010111000100111","001111011101001000110011010","001111011111010100010000010","001111100000010000010011110","001111100000101101110100000","001111100000100000110000010","001111100000001101111011000","001111011111011011111000011","001111011110001111011111011","001111011011010101111011110","001111011010000100011001000","001111011001101001110000000","001111011000011111101001010","001111011001100000010011100","001111011010000011110000000","000000000000000000000000000","000000000000000000000000000"),
                        ("000000000000000000000000000","001111011001100001111111100","001111011000000001110010110","001111010000111101101010110","001111001010010010110101010","001110111001110011101101000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","001111010001000011111011011","001111011001001010110111011","001111011100101001000011101","001111011100111101001111100","001111011001111111011101011","001111011000111001100010000","001111010011010001101110110","001111010100100111001111010","001111010101011110110010000","001111010111000100011001010","001111010111011100111010111","001111011010101110010111111","001111011011000100110000110","001111011100100000001001110","001111011011010101100010100","000000000000000000000000000","000000000000000000000000000"),
                        ("000000000000000000000000000","001111011011011001000000111","001111011010110010101001101","001111010100110011001001101","001111001101010010100111111","001111000011010010100010001","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","001110110101110111010110111","001111010110011110100100000","001111011011110110101101011","001111011110011100000100101","001111011111100100101100000","001111011101000100101000011","001111011010010011110101110","001111011000101010101111101","001111010111101001000110000","001111011001001101010011101","001111011001100000110001011","001111011010111001111000000","001111011101100101110011010","001111011111001110011000111","001111100000100111101110110","001111011101001110110011001","000000000000000000000000000","000000000000000000000000000"),
                        ("000000000000000000000000000","001111011010011101010101011","001111011100101101111000100","001111100000000000110101011","001111011111100001101000111","001111011111101101111011111","001111011110100101010101101","001111011101000100001111010","001111011100101001100110010","001111011101110000101000011","001111011110110101000010001","001111100000011100111101100","001111100001100100100100011","001111100011010101011001001","001111100100111100000101001","001111100101001111111010101","001111100100100101010110011","001111100001101010010101100","001111011100111011001101100","001111010100001011010110101","001110101010101011001001011","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","001111010101010110011110011","001111010010111101100111001","000000000000000000000000000","000000000000000000000000000"),
                        ("000000000000000000000000000","001111000100000001101001111","001110110010010101111010011","001111000011000011000100010","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","001110111001011011101101111","001111001110110101101101110","001111010011011000110011110","001111010011011110101010001","001111010010110000111110101","001111010010110011101010101","001111010000010110010111010","001111001110101001101100000","001111001111110000111111100","001111001101111010111001010","001111010001011001001110100","001111010010110001100100011","001111010101010001101000000","001111011000011000100010110","001111011001000110010011111","001111010001100111110000101","000000000000000000000000000","000000000000000000000000000"),
                        ("000000000000000000000000000","001111010111101100110100000","001111011100100010001001001","001111011110101110000010011","001111011110011000011001010","001111011101011010101101011","001111011100101011010111000","001111011101101100000110100","001111011110110101101000100","001111011110110010101100010","001111011110101110000100100","001111011110011011000110010","001111011110011101111100010","001111011110011111000100000","001111011101001010011001000","001111011100000011010101111","001111011010000000000101110","001111011000111100100001011","001111010011110111000011011","001111000100000100101111000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","001111000011001010001101100","001111011001100011000011101","000000000000000000000000000","000000000000000000000000000"),
                        ("000000000000000000000000000","001111001011010011000001101","001111001111111111101101001","001111000000110111100010101","001111001000001111101110101","001111010000001010000000101","001111010010101000000000000","001111010100100101000011111","001111010010010000001001010","001111010001011010000101000","001111010000000100111111110","001111001100110000101111100","001111000101001101110011101","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000"),
                        ("000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000"),
                        ("000000000000000000000000000","001111010110111111010010000","001111011011010100000100110","001111011110100100010010100","001111011110111000110001110","001111011111001101101111011","001111011111000101001010000","001111011110111100101111100","001111011111101001010000100","001111100000000010001010101","001111011111111110110111000","001111100000000111111101010","001111011111010110110010010","001111011111011000110110011","001111011110011011100001100","001111011100101110000011000","001111011001111100100101111","001111010011111101011100011","001111001011110011011001101","001111000010011010000010101","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","001111000010011011000001101","001111001110111100011011101","001111011000000001010101011","001111011000110001101110011","001111011010110010001001101","001111011100111000110010010","001111100000010110010101101","000000000000000000000000000","000000000000000000000000000"),
                        ("000000000000000000000000000","001111100001010010101111110","001111100011000010111101110","001111100010110101110000111","001111100011000000101101100","001111100010101000010010001","001111100010110010110110110","001111100010011010011001100","001111100001111101011010100","001111100001000001011011011","001111011110101100011000000","001111011101101110001100001","001111011100000100110010001","001111011011010010110001111","001111011011100000001011001","001111011101010001110011000","001111100001000010101111111","001111100100001000011111001","001111100101000101111001011","001111100111011001011011101","001111101000011010100101001","001111101001010010111101110","001111101001111000000000111","001111101010011001000010011","001111101010010100100000110","001111101010000111001110100","001111101001101010110111000","001111101000110111100100100","001111101000101010001111000","001111100101000111110000001","000000000000000000000000000","000000000000000000000000000"),
                        ("000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","001111001101111011011000110","001111011011110000111001101","001111100001100001000000100","001111100100011000001010001","001111100111110101101011011","001111101001011111000010111","001111101010100000011110010","001111101010111000111110011","001111101010010001110101010","001111101000110101001110101","001111100110100111110011100","001111100011011010000010011","001111011111101101001010101","001111010010100011110110110","000000000000000000000000000","000000000000000000000000000"),
                        ("000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","001111000001110111100100100","001111001110110000111001011","001111010110111101000001011","001111011010100100111101100","001111011111111101001011101","001111100001010011010100000","001111100010110111001100011","001111100001111110111110101","001111100010000001100001110","001111011111100000110011100","001111011011100001111011010","001111011000100010110101110","001111001100011111111011101","001111000101110111101011110","000000000000000000000000000","000000000000000000000000000"),
                        ("000000000000000000000000000","001111100001001010001011101","001111100100101001100011001","001111100101110101100011100","001111100101011111110001011","001111100101001010011110110","001111100101010000011111011","001111100100011001010111011","001111100100011100111001001","001111100011111011101101000","001111100011100111101011011","001111100011110111111000001","001111100100010000100111010","001111100100011110100000101","001111100101011011111011100","001111100101001111000010000","001111100100011010110110010","001111100010111001111101010","001111100001011001110000111","001111011111001101001001001","001111011101010100010001010","001111011010010011111100101","001111011011011110111000110","001111011111001101100111101","001111100000101110011011101","001111100010110010001101111","001111100011111011001011111","001111100101110010110010000","001111100110101110101011111","001111100110011100110101001","000000000000000000000000000","000000000000000000000000000"),
                        ("000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000"),
                        ("000000000000000000000000000","001111010011111100011101100","001111001000001000111100100","001111000111011111101100001","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","001111001011111101011111100","001111011010010100110100101","001111100000001010000111110","001111100011100111100111011","001111100110111011000000001","001111101000010001000110011","001111101001100111110100000","001111101010110010001100010","001111101011011100011111000","001111101011010100001110011","001111101011000011110100001","001111101010000100100110100","001111101000111011101111001","001111100111101000100000000","001111100101011011100001110","001111100001110110000011010","000000000000000000000000000","000000000000000000000000000"),
                        ("000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","001110110101000001111000010","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000"),
                        ("000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000"),
                        ("000000000000000000000000000","001111001111110101000101101","001111011000001001000111000","001111010000000000100101101","001111001000001011100100010","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","001111010000000011100100100","001111010010011111110001101","001111010010011100100111010","001111010010110111000101110","001111001101001011111110001","001110110101011111001111010","000000000000000000000000000","001110110100101000001100001","001111001110001000110010100","001111010110000111011110101","001111011000010111010111010","001111011011011010001000001","001111011110001010100001101","001111011111010011101100001","001111100000010101010100101","000000000000000000000000000","000000000000000000000000000"),
                        ("000000000000000000000000000","001111010101101000011000011","001111010111010101011101111","001111011010000011101011011","001111011100011111110001101","001111011100100000011000100","001111011100111001010100011","001111011101111101100010101","001111011111010011101100001","001111100000011001001000010","001111100001000101000010101","001111100001101110111111010","001111100010100000101111110","001111100011001001000111100","001111100010111110010100110","001111100010100100001110101","001111100001011100000101100","001111100000010001001010011","001111011110000000100001000","001111011100101010110100111","001111011100011010111011110","001111011011101100000111100","001111011010110000111100100","001111011000010000011010001","001111011000010100100111101","001111010101000011010100100","001111010101001010000100100","001111010111011010111011000","001111010100000111011001111","001111010111000101000101010","000000000000000000000000000","000000000000000000000000000"),
                        ("000000000000000000000000000","001111010010000111111101000","001111001111111100101100001","001111010000010000000100101","001111001000011001010011000","001110111011111101110110101","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","001111000100011001101101001","001111010010111010010000001","001111011010010000101001111","001111011110011100111111111","001111011110111101100101000","001111100000100001011001100","001111100000000111000001000","001111100000010001111011011","001111100000000000100101011","001111100000100000111110100","001111011111111010001010101","001111011111110100001000010","001111011111010101000101110","001111011110111011000110101","001111011111011001010011010","001111011110010110001011001","001111011011100000011001010","000000000000000000000000000","000000000000000000000000000"),
                        ("000000000000000000000000000","001111100010101100011011101","001111100011011000111110010","001111100100001011011101011","001111100011110111001110001","001111100011110110100111001","001111100100000101011110011","001111100011101111101011010","001111100011000000110011111","001111100001111001111111101","001111100010001111001001111","001111100010001000011001011","001111100001110111100101000","001111100010000000100111110","001111100010011100110001000","001111100010111010111101010","001111100010110001011011000","001111011111111001110000011","001111011101100011101101000","001111010111010111100011000","001111010000001110011001101","001111000001000101001011000","001111001010011011000001101","001111001001001011101110100","001111010101100010010010011","001111011010011100110010010","001111011101011010110010001","001111100001100010100010111","001111100010100000110001101","001111100010001001111011011","000000000000000000000000000","000000000000000000000000000"),
                        ("000000000000000000000000000","001110111100110100100000101","001111001000110010111101000","001111010010111100101011011","001111010011110001101010011","001111010100010011000001011","001111010110100101011011011","001111011000001011100110011","001111011001010101101011100","001111011001101000110010001","001111011000100001110111111","001111010110010001011010000","001111010000101111110111111","001111001000111101000000111","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000"),
                        ("000000000000000000000000000","001111100001000101101100101","001111100000111000000000100","001111100001011111011100101","001111100001000101010101100","001111100001001010010011100","001111100001000011001100101","001111100001000101101100111","001111100000101010111110011","001111011111101011110001000","001111011110010110110110110","001111011100101011110010010","001111011011111001000001010","001111011010100111010000011","001111011010011011010101100","001111011100000111011001011","001111011101100110101110000","001111011101100110110011110","001111011100001111010001010","001111011001000101001110110","001111010101010101111010101","001111001111110010011111111","001111001100011011000101010","001111001111000000011001011","001111010101110110011110010","001111011000110001001000001","001111011011111011001100110","001111011110100100101101110","001111100000100011110000110","001111011100101001110011111","000000000000000000000000000","000000000000000000000000000"),
                        ("000000000000000000000000000","001111100010001000101110010","001111100011001100011000101","001111100011100001000101000","001111100010101000010001011","001111100010011011010100110","001111100010010111000111010","001111100010011011100101000","001111100010010111000001100","001111100001111101100100100","001111100000101001111000101","001111011110000011010001101","001111011011010001000110111","001111011000100001101111100","001111010001101101111111000","001111001000010100101101011","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","000000000000000000000000000","001111001110001110100111110","001111011001001000010000001","001111011101110101111100101","001111100000100101001110000","001111100001110110011100101","001111011111110110001011011","000000000000000000000000000","000000000000000000000000000"));    
      
        wait for 300ns;
        wait;
        
    end process;
         

end Behavioral;
